

module image_cell (
 input clk, 
 input GlobalReset, 
 input Input_Valid,
 //input valid_max, //
 input [9:0] Pix_0, // sfix10_En0 
 input [9:0] Pix_1, // sfix10_En0 
 input [9:0] Pix_2, // sfix10_En0 
 input [9:0] Pix_3, // sfix10_En0 
 input [9:0] Pix_4, // sfix10_En0 
 input [9:0] Pix_5, // sfix10_En0 
 input [9:0] Pix_6, // sfix10_En0 
 input [9:0] Pix_7, // sfix10_En0 
 input [9:0] Pix_8, // sfix10_En0 
 input [9:0] Pix_9, // sfix10_En0 
 input [9:0] Pix_10, // sfix10_En0 
 input [9:0] Pix_11, // sfix10_En0 
 input [9:0] Pix_12, // sfix10_En0 
 input [9:0] Pix_13, // sfix10_En0 
 input [9:0] Pix_14, // sfix10_En0 
 input [9:0] Pix_15, // sfix10_En0 
 input [9:0] Pix_16, // sfix10_En0 
 input [9:0] Pix_17, // sfix10_En0 
 input [9:0] Pix_18, // sfix10_En0 
 input [9:0] Pix_19, // sfix10_En0 
 input [9:0] Pix_20, // sfix10_En0 
 input [9:0] Pix_21, // sfix10_En0 
 input [9:0] Pix_22, // sfix10_En0 
 input [9:0] Pix_23, // sfix10_En0 
 input [9:0] Pix_24, // sfix10_En0 
 input [9:0] Pix_25, // sfix10_En0 
 input [9:0] Pix_26, // sfix10_En0 
 input [9:0] Pix_27, // sfix10_En0 
 input [9:0] Pix_28, // sfix10_En0 
 input [9:0] Pix_29, // sfix10_En0 
 input [9:0] Pix_30, // sfix10_En0 
 input [9:0] Pix_31, // sfix10_En0 
 input [9:0] Pix_32, // sfix10_En0 
 input [9:0] Pix_33, // sfix10_En0 
 input [9:0] Pix_34, // sfix10_En0 
 input [9:0] Pix_35, // sfix10_En0 
 input [9:0] Pix_36, // sfix10_En0 
 input [9:0] Pix_37, // sfix10_En0 
 input [9:0] Pix_38, // sfix10_En0 
 input [9:0] Pix_39, // sfix10_En0 
 input [9:0] Pix_40, // sfix10_En0 
 input [9:0] Pix_41, // sfix10_En0 
 input [9:0] Pix_42, // sfix10_En0 
 input [9:0] Pix_43, // sfix10_En0 
 input [9:0] Pix_44, // sfix10_En0 
 input [9:0] Pix_45, // sfix10_En0 
 input [9:0] Pix_46, // sfix10_En0 
 input [9:0] Pix_47, // sfix10_En0 
 input [9:0] Pix_48, // sfix10_En0 
 input [9:0] Pix_49, // sfix10_En0 
 input [9:0] Pix_50, // sfix10_En0 
 input [9:0] Pix_51, // sfix10_En0 
 input [9:0] Pix_52, // sfix10_En0 
 input [9:0] Pix_53, // sfix10_En0 
 input [9:0] Pix_54, // sfix10_En0 
 input [9:0] Pix_55, // sfix10_En0 
 input [9:0] Pix_56, // sfix10_En0 
 input [9:0] Pix_57, // sfix10_En0 
 input [9:0] Pix_58, // sfix10_En0 
 input [9:0] Pix_59, // sfix10_En0 
 input [9:0] Pix_60, // sfix10_En0 
 input [9:0] Pix_61, // sfix10_En0 
 input [9:0] Pix_62, // sfix10_En0 
 input [9:0] Pix_63, // sfix10_En0 
 input [9:0] Pix_64, // sfix10_En0 
 input [9:0] Pix_65, // sfix10_En0 
 input [9:0] Pix_66, // sfix10_En0 
 input [9:0] Pix_67, // sfix10_En0 
 input [9:0] Pix_68, // sfix10_En0 
 input [9:0] Pix_69, // sfix10_En0 
 input [9:0] Pix_70, // sfix10_En0 
 input [9:0] Pix_71, // sfix10_En0 
 input [9:0] Pix_72, // sfix10_En0 
 input [9:0] Pix_73, // sfix10_En0 
 input [9:0] Pix_74, // sfix10_En0 
 input [9:0] Pix_75, // sfix10_En0 
 input [9:0] Pix_76, // sfix10_En0 
 input [9:0] Pix_77, // sfix10_En0 
 input [9:0] Pix_78, // sfix10_En0 
 input [9:0] Pix_79, // sfix10_En0 
 input [9:0] Pix_80, // sfix10_En0 
 input [9:0] Pix_81, // sfix10_En0 
 input [9:0] Pix_82, // sfix10_En0 
 input [9:0] Pix_83, // sfix10_En0 
 input [9:0] Pix_84, // sfix10_En0 
 input [9:0] Pix_85, // sfix10_En0 
 input [9:0] Pix_86, // sfix10_En0 
 input [9:0] Pix_87, // sfix10_En0 
 input [9:0] Pix_88, // sfix10_En0 
 input [9:0] Pix_89, // sfix10_En0 
 input [9:0] Pix_90, // sfix10_En0 
 input [9:0] Pix_91, // sfix10_En0 
 input [9:0] Pix_92, // sfix10_En0 
 input [9:0] Pix_93, // sfix10_En0 
 input [9:0] Pix_94, // sfix10_En0 
 input [9:0] Pix_95, // sfix10_En0 
 input [9:0] Pix_96, // sfix10_En0 
 input [9:0] Pix_97, // sfix10_En0 
 input [9:0] Pix_98, // sfix10_En0 
 input [9:0] Pix_99, // sfix10_En0 
 input [9:0] Pix_100, // sfix10_En0 
 input [9:0] Pix_101, // sfix10_En0 
 input [9:0] Pix_102, // sfix10_En0 
 input [9:0] Pix_103, // sfix10_En0 
 input [9:0] Pix_104, // sfix10_En0 
 input [9:0] Pix_105, // sfix10_En0 
 input [9:0] Pix_106, // sfix10_En0 
 input [9:0] Pix_107, // sfix10_En0 
 input [9:0] Pix_108, // sfix10_En0 
 input [9:0] Pix_109, // sfix10_En0 
 input [9:0] Pix_110, // sfix10_En0 
 input [9:0] Pix_111, // sfix10_En0 
 input [9:0] Pix_112, // sfix10_En0 
 input [9:0] Pix_113, // sfix10_En0 
 input [9:0] Pix_114, // sfix10_En0 
 input [9:0] Pix_115, // sfix10_En0 
 input [9:0] Pix_116, // sfix10_En0 
 input [9:0] Pix_117, // sfix10_En0 
 input [9:0] Pix_118, // sfix10_En0 
 input [9:0] Pix_119, // sfix10_En0 
 input [9:0] Pix_120, // sfix10_En0 
 input [9:0] Pix_121, // sfix10_En0 
 input [9:0] Pix_122, // sfix10_En0 
 input [9:0] Pix_123, // sfix10_En0 
 input [9:0] Pix_124, // sfix10_En0 
 input [9:0] Pix_125, // sfix10_En0 
 input [9:0] Pix_126, // sfix10_En0 
 input [9:0] Pix_127, // sfix10_En0 
 input [9:0] Pix_128, // sfix10_En0 
 input [9:0] Pix_129, // sfix10_En0 
 input [9:0] Pix_130, // sfix10_En0 
 input [9:0] Pix_131, // sfix10_En0 
 input [9:0] Pix_132, // sfix10_En0 
 input [9:0] Pix_133, // sfix10_En0 
 input [9:0] Pix_134, // sfix10_En0 
 input [9:0] Pix_135, // sfix10_En0 
 input [9:0] Pix_136, // sfix10_En0 
 input [9:0] Pix_137, // sfix10_En0 
 input [9:0] Pix_138, // sfix10_En0 
 input [9:0] Pix_139, // sfix10_En0 
 input [9:0] Pix_140, // sfix10_En0 
 input [9:0] Pix_141, // sfix10_En0 
 input [9:0] Pix_142, // sfix10_En0 
 input [9:0] Pix_143, // sfix10_En0 
 input [9:0] Pix_144, // sfix10_En0 
 input [9:0] Pix_145, // sfix10_En0 
 input [9:0] Pix_146, // sfix10_En0 
 input [9:0] Pix_147, // sfix10_En0 
 input [9:0] Pix_148, // sfix10_En0 
 input [9:0] Pix_149, // sfix10_En0 
 input [9:0] Pix_150, // sfix10_En0 
 input [9:0] Pix_151, // sfix10_En0 
 input [9:0] Pix_152, // sfix10_En0 
 input [9:0] Pix_153, // sfix10_En0 
 input [9:0] Pix_154, // sfix10_En0 
 input [9:0] Pix_155, // sfix10_En0 
 input [9:0] Pix_156, // sfix10_En0 
 input [9:0] Pix_157, // sfix10_En0 
 input [9:0] Pix_158, // sfix10_En0 
 input [9:0] Pix_159, // sfix10_En0 
 input [9:0] Pix_160, // sfix10_En0 
 input [9:0] Pix_161, // sfix10_En0 
 input [9:0] Pix_162, // sfix10_En0 
 input [9:0] Pix_163, // sfix10_En0 
 input [9:0] Pix_164, // sfix10_En0 
 input [9:0] Pix_165, // sfix10_En0 
 input [9:0] Pix_166, // sfix10_En0 
 input [9:0] Pix_167, // sfix10_En0 
 input [9:0] Pix_168, // sfix10_En0 
 input [9:0] Pix_169, // sfix10_En0 
 input [9:0] Pix_170, // sfix10_En0 
 input [9:0] Pix_171, // sfix10_En0 
 input [9:0] Pix_172, // sfix10_En0 
 input [9:0] Pix_173, // sfix10_En0 
 input [9:0] Pix_174, // sfix10_En0 
 input [9:0] Pix_175, // sfix10_En0 
 input [9:0] Pix_176, // sfix10_En0 
 input [9:0] Pix_177, // sfix10_En0 
 input [9:0] Pix_178, // sfix10_En0 
 input [9:0] Pix_179, // sfix10_En0 
 input [9:0] Pix_180, // sfix10_En0 
 input [9:0] Pix_181, // sfix10_En0 
 input [9:0] Pix_182, // sfix10_En0 
 input [9:0] Pix_183, // sfix10_En0 
 input [9:0] Pix_184, // sfix10_En0 
 input [9:0] Pix_185, // sfix10_En0 
 input [9:0] Pix_186, // sfix10_En0 
 input [9:0] Pix_187, // sfix10_En0 
 input [9:0] Pix_188, // sfix10_En0 
 input [9:0] Pix_189, // sfix10_En0 
 input [9:0] Pix_190, // sfix10_En0 
 input [9:0] Pix_191, // sfix10_En0 
 input [9:0] Pix_192, // sfix10_En0 
 input [9:0] Pix_193, // sfix10_En0 
 input [9:0] Pix_194, // sfix10_En0 
 input [9:0] Pix_195, // sfix10_En0 
 input [9:0] Pix_196, // sfix10_En0 
 input [9:0] Pix_197, // sfix10_En0 
 input [9:0] Pix_198, // sfix10_En0 
 input [9:0] Pix_199, // sfix10_En0 
 input [9:0] Pix_200, // sfix10_En0 
 input [9:0] Pix_201, // sfix10_En0 
 input [9:0] Pix_202, // sfix10_En0 
 input [9:0] Pix_203, // sfix10_En0 
 input [9:0] Pix_204, // sfix10_En0 
 input [9:0] Pix_205, // sfix10_En0 
 input [9:0] Pix_206, // sfix10_En0 
 input [9:0] Pix_207, // sfix10_En0 
 input [9:0] Pix_208, // sfix10_En0 
 input [9:0] Pix_209, // sfix10_En0 
 input [9:0] Pix_210, // sfix10_En0 
 input [9:0] Pix_211, // sfix10_En0 
 input [9:0] Pix_212, // sfix10_En0 
 input [9:0] Pix_213, // sfix10_En0 
 input [9:0] Pix_214, // sfix10_En0 
 input [9:0] Pix_215, // sfix10_En0 
 input [9:0] Pix_216, // sfix10_En0 
 input [9:0] Pix_217, // sfix10_En0 
 input [9:0] Pix_218, // sfix10_En0 
 input [9:0] Pix_219, // sfix10_En0 
 input [9:0] Pix_220, // sfix10_En0 
 input [9:0] Pix_221, // sfix10_En0 
 input [9:0] Pix_222, // sfix10_En0 
 input [9:0] Pix_223, // sfix10_En0 
 input [9:0] Pix_224, // sfix10_En0 
 input [9:0] Pix_225, // sfix10_En0 
 input [9:0] Pix_226, // sfix10_En0 
 input [9:0] Pix_227, // sfix10_En0 
 input [9:0] Pix_228, // sfix10_En0 
 input [9:0] Pix_229, // sfix10_En0 
 input [9:0] Pix_230, // sfix10_En0 
 input [9:0] Pix_231, // sfix10_En0 
 input [9:0] Pix_232, // sfix10_En0 
 input [9:0] Pix_233, // sfix10_En0 
 input [9:0] Pix_234, // sfix10_En0 
 input [9:0] Pix_235, // sfix10_En0 
 input [9:0] Pix_236, // sfix10_En0 
 input [9:0] Pix_237, // sfix10_En0 
 input [9:0] Pix_238, // sfix10_En0 
 input [9:0] Pix_239, // sfix10_En0 
 input [9:0] Pix_240, // sfix10_En0 
 input [9:0] Pix_241, // sfix10_En0 
 input [9:0] Pix_242, // sfix10_En0 
 input [9:0] Pix_243, // sfix10_En0 
 input [9:0] Pix_244, // sfix10_En0 
 input [9:0] Pix_245, // sfix10_En0 
 input [9:0] Pix_246, // sfix10_En0 
 input [9:0] Pix_247, // sfix10_En0 
 input [9:0] Pix_248, // sfix10_En0 
 input [9:0] Pix_249, // sfix10_En0 
 input [9:0] Pix_250, // sfix10_En0 
 input [9:0] Pix_251, // sfix10_En0 
 input [9:0] Pix_252, // sfix10_En0 
 input [9:0] Pix_253, // sfix10_En0 
 input [9:0] Pix_254, // sfix10_En0 
 input [9:0] Pix_255, // sfix10_En0 
 input [9:0] Pix_256, // sfix10_En0 
 input [9:0] Pix_257, // sfix10_En0 
 input [9:0] Pix_258, // sfix10_En0 
 input [9:0] Pix_259, // sfix10_En0 
 input [9:0] Pix_260, // sfix10_En0 
 input [9:0] Pix_261, // sfix10_En0 
 input [9:0] Pix_262, // sfix10_En0 
 input [9:0] Pix_263, // sfix10_En0 
 input [9:0] Pix_264, // sfix10_En0 
 input [9:0] Pix_265, // sfix10_En0 
 input [9:0] Pix_266, // sfix10_En0 
 input [9:0] Pix_267, // sfix10_En0 
 input [9:0] Pix_268, // sfix10_En0 
 input [9:0] Pix_269, // sfix10_En0 
 input [9:0] Pix_270, // sfix10_En0 
 input [9:0] Pix_271, // sfix10_En0 
 input [9:0] Pix_272, // sfix10_En0 
 input [9:0] Pix_273, // sfix10_En0 
 input [9:0] Pix_274, // sfix10_En0 
 input [9:0] Pix_275, // sfix10_En0 
 input [9:0] Pix_276, // sfix10_En0 
 input [9:0] Pix_277, // sfix10_En0 
 input [9:0] Pix_278, // sfix10_En0 
 input [9:0] Pix_279, // sfix10_En0 
 input [9:0] Pix_280, // sfix10_En0 
 input [9:0] Pix_281, // sfix10_En0 
 input [9:0] Pix_282, // sfix10_En0 
 input [9:0] Pix_283, // sfix10_En0 
 input [9:0] Pix_284, // sfix10_En0 
 input [9:0] Pix_285, // sfix10_En0 
 input [9:0] Pix_286, // sfix10_En0 
 input [9:0] Pix_287, // sfix10_En0 
 input [9:0] Pix_288, // sfix10_En0 
 input [9:0] Pix_289, // sfix10_En0 
 input [9:0] Pix_290, // sfix10_En0 
 input [9:0] Pix_291, // sfix10_En0 
 input [9:0] Pix_292, // sfix10_En0 
 input [9:0] Pix_293, // sfix10_En0 
 input [9:0] Pix_294, // sfix10_En0 
 input [9:0] Pix_295, // sfix10_En0 
 input [9:0] Pix_296, // sfix10_En0 
 input [9:0] Pix_297, // sfix10_En0 
 input [9:0] Pix_298, // sfix10_En0 
 input [9:0] Pix_299, // sfix10_En0 
 input [9:0] Pix_300, // sfix10_En0 
 input [9:0] Pix_301, // sfix10_En0 
 input [9:0] Pix_302, // sfix10_En0 
 input [9:0] Pix_303, // sfix10_En0 
 input [9:0] Pix_304, // sfix10_En0 
 input [9:0] Pix_305, // sfix10_En0 
 input [9:0] Pix_306, // sfix10_En0 
 input [9:0] Pix_307, // sfix10_En0 
 input [9:0] Pix_308, // sfix10_En0 
 input [9:0] Pix_309, // sfix10_En0 
 input [9:0] Pix_310, // sfix10_En0 
 input [9:0] Pix_311, // sfix10_En0 
 input [9:0] Pix_312, // sfix10_En0 
 input [9:0] Pix_313, // sfix10_En0 
 input [9:0] Pix_314, // sfix10_En0 
 input [9:0] Pix_315, // sfix10_En0 
 input [9:0] Pix_316, // sfix10_En0 
 input [9:0] Pix_317, // sfix10_En0 
 input [9:0] Pix_318, // sfix10_En0 
 input [9:0] Pix_319, // sfix10_En0 
 input [9:0] Pix_320, // sfix10_En0 
 input [9:0] Pix_321, // sfix10_En0 
 input [9:0] Pix_322, // sfix10_En0 
 input [9:0] Pix_323, // sfix10_En0 
 input [9:0] Pix_324, // sfix10_En0 
 input [9:0] Pix_325, // sfix10_En0 
 input [9:0] Pix_326, // sfix10_En0 
 input [9:0] Pix_327, // sfix10_En0 
 input [9:0] Pix_328, // sfix10_En0 
 input [9:0] Pix_329, // sfix10_En0 
 input [9:0] Pix_330, // sfix10_En0 
 input [9:0] Pix_331, // sfix10_En0 
 input [9:0] Pix_332, // sfix10_En0 
 input [9:0] Pix_333, // sfix10_En0 
 input [9:0] Pix_334, // sfix10_En0 
 input [9:0] Pix_335, // sfix10_En0 
 input [9:0] Pix_336, // sfix10_En0 
 input [9:0] Pix_337, // sfix10_En0 
 input [9:0] Pix_338, // sfix10_En0 
 input [9:0] Pix_339, // sfix10_En0 
 input [9:0] Pix_340, // sfix10_En0 
 input [9:0] Pix_341, // sfix10_En0 
 input [9:0] Pix_342, // sfix10_En0 
 input [9:0] Pix_343, // sfix10_En0 
 input [9:0] Pix_344, // sfix10_En0 
 input [9:0] Pix_345, // sfix10_En0 
 input [9:0] Pix_346, // sfix10_En0 
 input [9:0] Pix_347, // sfix10_En0 
 input [9:0] Pix_348, // sfix10_En0 
 input [9:0] Pix_349, // sfix10_En0 
 input [9:0] Pix_350, // sfix10_En0 
 input [9:0] Pix_351, // sfix10_En0 
 input [9:0] Pix_352, // sfix10_En0 
 input [9:0] Pix_353, // sfix10_En0 
 input [9:0] Pix_354, // sfix10_En0 
 input [9:0] Pix_355, // sfix10_En0 
 input [9:0] Pix_356, // sfix10_En0 
 input [9:0] Pix_357, // sfix10_En0 
 input [9:0] Pix_358, // sfix10_En0 
 input [9:0] Pix_359, // sfix10_En0 
 input [9:0] Pix_360, // sfix10_En0 
 input [9:0] Pix_361, // sfix10_En0 
 input [9:0] Pix_362, // sfix10_En0 
 input [9:0] Pix_363, // sfix10_En0 
 input [9:0] Pix_364, // sfix10_En0 
 input [9:0] Pix_365, // sfix10_En0 
 input [9:0] Pix_366, // sfix10_En0 
 input [9:0] Pix_367, // sfix10_En0 
 input [9:0] Pix_368, // sfix10_En0 
 input [9:0] Pix_369, // sfix10_En0 
 input [9:0] Pix_370, // sfix10_En0 
 input [9:0] Pix_371, // sfix10_En0 
 input [9:0] Pix_372, // sfix10_En0 
 input [9:0] Pix_373, // sfix10_En0 
 input [9:0] Pix_374, // sfix10_En0 
 input [9:0] Pix_375, // sfix10_En0 
 input [9:0] Pix_376, // sfix10_En0 
 input [9:0] Pix_377, // sfix10_En0 
 input [9:0] Pix_378, // sfix10_En0 
 input [9:0] Pix_379, // sfix10_En0 
 input [9:0] Pix_380, // sfix10_En0 
 input [9:0] Pix_381, // sfix10_En0 
 input [9:0] Pix_382, // sfix10_En0 
 input [9:0] Pix_383, // sfix10_En0 
 input [9:0] Pix_384, // sfix10_En0 
 input [9:0] Pix_385, // sfix10_En0 
 input [9:0] Pix_386, // sfix10_En0 
 input [9:0] Pix_387, // sfix10_En0 
 input [9:0] Pix_388, // sfix10_En0 
 input [9:0] Pix_389, // sfix10_En0 
 input [9:0] Pix_390, // sfix10_En0 
 input [9:0] Pix_391, // sfix10_En0 
 input [9:0] Pix_392, // sfix10_En0 
 input [9:0] Pix_393, // sfix10_En0 
 input [9:0] Pix_394, // sfix10_En0 
 input [9:0] Pix_395, // sfix10_En0 
 input [9:0] Pix_396, // sfix10_En0 
 input [9:0] Pix_397, // sfix10_En0 
 input [9:0] Pix_398, // sfix10_En0 
 input [9:0] Pix_399, // sfix10_En0 
 input [9:0] Pix_400, // sfix10_En0 
 input [9:0] Pix_401, // sfix10_En0 
 input [9:0] Pix_402, // sfix10_En0 
 input [9:0] Pix_403, // sfix10_En0 
 input [9:0] Pix_404, // sfix10_En0 
 input [9:0] Pix_405, // sfix10_En0 
 input [9:0] Pix_406, // sfix10_En0 
 input [9:0] Pix_407, // sfix10_En0 
 input [9:0] Pix_408, // sfix10_En0 
 input [9:0] Pix_409, // sfix10_En0 
 input [9:0] Pix_410, // sfix10_En0 
 input [9:0] Pix_411, // sfix10_En0 
 input [9:0] Pix_412, // sfix10_En0 
 input [9:0] Pix_413, // sfix10_En0 
 input [9:0] Pix_414, // sfix10_En0 
 input [9:0] Pix_415, // sfix10_En0 
 input [9:0] Pix_416, // sfix10_En0 
 input [9:0] Pix_417, // sfix10_En0 
 input [9:0] Pix_418, // sfix10_En0 
 input [9:0] Pix_419, // sfix10_En0 
 input [9:0] Pix_420, // sfix10_En0 
 input [9:0] Pix_421, // sfix10_En0 
 input [9:0] Pix_422, // sfix10_En0 
 input [9:0] Pix_423, // sfix10_En0 
 input [9:0] Pix_424, // sfix10_En0 
 input [9:0] Pix_425, // sfix10_En0 
 input [9:0] Pix_426, // sfix10_En0 
 input [9:0] Pix_427, // sfix10_En0 
 input [9:0] Pix_428, // sfix10_En0 
 input [9:0] Pix_429, // sfix10_En0 
 input [9:0] Pix_430, // sfix10_En0 
 input [9:0] Pix_431, // sfix10_En0 
 input [9:0] Pix_432, // sfix10_En0 
 input [9:0] Pix_433, // sfix10_En0 
 input [9:0] Pix_434, // sfix10_En0 
 input [9:0] Pix_435, // sfix10_En0 
 input [9:0] Pix_436, // sfix10_En0 
 input [9:0] Pix_437, // sfix10_En0 
 input [9:0] Pix_438, // sfix10_En0 
 input [9:0] Pix_439, // sfix10_En0 
 input [9:0] Pix_440, // sfix10_En0 
 input [9:0] Pix_441, // sfix10_En0 
 input [9:0] Pix_442, // sfix10_En0 
 input [9:0] Pix_443, // sfix10_En0 
 input [9:0] Pix_444, // sfix10_En0 
 input [9:0] Pix_445, // sfix10_En0 
 input [9:0] Pix_446, // sfix10_En0 
 input [9:0] Pix_447, // sfix10_En0 
 input [9:0] Pix_448, // sfix10_En0 
 input [9:0] Pix_449, // sfix10_En0 
 input [9:0] Pix_450, // sfix10_En0 
 input [9:0] Pix_451, // sfix10_En0 
 input [9:0] Pix_452, // sfix10_En0 
 input [9:0] Pix_453, // sfix10_En0 
 input [9:0] Pix_454, // sfix10_En0 
 input [9:0] Pix_455, // sfix10_En0 
 input [9:0] Pix_456, // sfix10_En0 
 input [9:0] Pix_457, // sfix10_En0 
 input [9:0] Pix_458, // sfix10_En0 
 input [9:0] Pix_459, // sfix10_En0 
 input [9:0] Pix_460, // sfix10_En0 
 input [9:0] Pix_461, // sfix10_En0 
 input [9:0] Pix_462, // sfix10_En0 
 input [9:0] Pix_463, // sfix10_En0 
 input [9:0] Pix_464, // sfix10_En0 
 input [9:0] Pix_465, // sfix10_En0 
 input [9:0] Pix_466, // sfix10_En0 
 input [9:0] Pix_467, // sfix10_En0 
 input [9:0] Pix_468, // sfix10_En0 
 input [9:0] Pix_469, // sfix10_En0 
 input [9:0] Pix_470, // sfix10_En0 
 input [9:0] Pix_471, // sfix10_En0 
 input [9:0] Pix_472, // sfix10_En0 
 input [9:0] Pix_473, // sfix10_En0 
 input [9:0] Pix_474, // sfix10_En0 
 input [9:0] Pix_475, // sfix10_En0 
 input [9:0] Pix_476, // sfix10_En0 
 input [9:0] Pix_477, // sfix10_En0 
 input [9:0] Pix_478, // sfix10_En0 
 input [9:0] Pix_479, // sfix10_En0 
 input [9:0] Pix_480, // sfix10_En0 
 input [9:0] Pix_481, // sfix10_En0 
 input [9:0] Pix_482, // sfix10_En0 
 input [9:0] Pix_483, // sfix10_En0 
 input [9:0] Pix_484, // sfix10_En0 
 input [9:0] Pix_485, // sfix10_En0 
 input [9:0] Pix_486, // sfix10_En0 
 input [9:0] Pix_487, // sfix10_En0 
 input [9:0] Pix_488, // sfix10_En0 
 input [9:0] Pix_489, // sfix10_En0 
 input [9:0] Pix_490, // sfix10_En0 
 input [9:0] Pix_491, // sfix10_En0 
 input [9:0] Pix_492, // sfix10_En0 
 input [9:0] Pix_493, // sfix10_En0 
 input [9:0] Pix_494, // sfix10_En0 
 input [9:0] Pix_495, // sfix10_En0 
 input [9:0] Pix_496, // sfix10_En0 
 input [9:0] Pix_497, // sfix10_En0 
 input [9:0] Pix_498, // sfix10_En0 
 input [9:0] Pix_499, // sfix10_En0 
 input [9:0] Pix_500, // sfix10_En0 
 input [9:0] Pix_501, // sfix10_En0 
 input [9:0] Pix_502, // sfix10_En0 
 input [9:0] Pix_503, // sfix10_En0 
 input [9:0] Pix_504, // sfix10_En0 
 input [9:0] Pix_505, // sfix10_En0 
 input [9:0] Pix_506, // sfix10_En0 
 input [9:0] Pix_507, // sfix10_En0 
 input [9:0] Pix_508, // sfix10_En0 
 input [9:0] Pix_509, // sfix10_En0 
 input [9:0] Pix_510, // sfix10_En0 
 input [9:0] Pix_511, // sfix10_En0 
 input [9:0] Pix_512, // sfix10_En0 
 input [9:0] Pix_513, // sfix10_En0 
 input [9:0] Pix_514, // sfix10_En0 
 input [9:0] Pix_515, // sfix10_En0 
 input [9:0] Pix_516, // sfix10_En0 
 input [9:0] Pix_517, // sfix10_En0 
 input [9:0] Pix_518, // sfix10_En0 
 input [9:0] Pix_519, // sfix10_En0 
 input [9:0] Pix_520, // sfix10_En0 
 input [9:0] Pix_521, // sfix10_En0 
 input [9:0] Pix_522, // sfix10_En0 
 input [9:0] Pix_523, // sfix10_En0 
 input [9:0] Pix_524, // sfix10_En0 
 input [9:0] Pix_525, // sfix10_En0 
 input [9:0] Pix_526, // sfix10_En0 
 input [9:0] Pix_527, // sfix10_En0 
 input [9:0] Pix_528, // sfix10_En0 
 input [9:0] Pix_529, // sfix10_En0 
 input [9:0] Pix_530, // sfix10_En0 
 input [9:0] Pix_531, // sfix10_En0 
 input [9:0] Pix_532, // sfix10_En0 
 input [9:0] Pix_533, // sfix10_En0 
 input [9:0] Pix_534, // sfix10_En0 
 input [9:0] Pix_535, // sfix10_En0 
 input [9:0] Pix_536, // sfix10_En0 
 input [9:0] Pix_537, // sfix10_En0 
 input [9:0] Pix_538, // sfix10_En0 
 input [9:0] Pix_539, // sfix10_En0 
 input [9:0] Pix_540, // sfix10_En0 
 input [9:0] Pix_541, // sfix10_En0 
 input [9:0] Pix_542, // sfix10_En0 
 input [9:0] Pix_543, // sfix10_En0 
 input [9:0] Pix_544, // sfix10_En0 
 input [9:0] Pix_545, // sfix10_En0 
 input [9:0] Pix_546, // sfix10_En0 
 input [9:0] Pix_547, // sfix10_En0 
 input [9:0] Pix_548, // sfix10_En0 
 input [9:0] Pix_549, // sfix10_En0 
 input [9:0] Pix_550, // sfix10_En0 
 input [9:0] Pix_551, // sfix10_En0 
 input [9:0] Pix_552, // sfix10_En0 
 input [9:0] Pix_553, // sfix10_En0 
 input [9:0] Pix_554, // sfix10_En0 
 input [9:0] Pix_555, // sfix10_En0 
 input [9:0] Pix_556, // sfix10_En0 
 input [9:0] Pix_557, // sfix10_En0 
 input [9:0] Pix_558, // sfix10_En0 
 input [9:0] Pix_559, // sfix10_En0 
 input [9:0] Pix_560, // sfix10_En0 
 input [9:0] Pix_561, // sfix10_En0 
 input [9:0] Pix_562, // sfix10_En0 
 input [9:0] Pix_563, // sfix10_En0 
 input [9:0] Pix_564, // sfix10_En0 
 input [9:0] Pix_565, // sfix10_En0 
 input [9:0] Pix_566, // sfix10_En0 
 input [9:0] Pix_567, // sfix10_En0 
 input [9:0] Pix_568, // sfix10_En0 
 input [9:0] Pix_569, // sfix10_En0 
 input [9:0] Pix_570, // sfix10_En0 
 input [9:0] Pix_571, // sfix10_En0 
 input [9:0] Pix_572, // sfix10_En0 
 input [9:0] Pix_573, // sfix10_En0 
 input [9:0] Pix_574, // sfix10_En0 
 input [9:0] Pix_575, // sfix10_En0 
 input [9:0] Pix_576, // sfix10_En0 
 input [9:0] Pix_577, // sfix10_En0 
 input [9:0] Pix_578, // sfix10_En0 
 input [9:0] Pix_579, // sfix10_En0 
 input [9:0] Pix_580, // sfix10_En0 
 input [9:0] Pix_581, // sfix10_En0 
 input [9:0] Pix_582, // sfix10_En0 
 input [9:0] Pix_583, // sfix10_En0 
 input [9:0] Pix_584, // sfix10_En0 
 input [9:0] Pix_585, // sfix10_En0 
 input [9:0] Pix_586, // sfix10_En0 
 input [9:0] Pix_587, // sfix10_En0 
 input [9:0] Pix_588, // sfix10_En0 
 input [9:0] Pix_589, // sfix10_En0 
 input [9:0] Pix_590, // sfix10_En0 
 input [9:0] Pix_591, // sfix10_En0 
 input [9:0] Pix_592, // sfix10_En0 
 input [9:0] Pix_593, // sfix10_En0 
 input [9:0] Pix_594, // sfix10_En0 
 input [9:0] Pix_595, // sfix10_En0 
 input [9:0] Pix_596, // sfix10_En0 
 input [9:0] Pix_597, // sfix10_En0 
 input [9:0] Pix_598, // sfix10_En0 
 input [9:0] Pix_599, // sfix10_En0 
 input [9:0] Pix_600, // sfix10_En0 
 input [9:0] Pix_601, // sfix10_En0 
 input [9:0] Pix_602, // sfix10_En0 
 input [9:0] Pix_603, // sfix10_En0 
 input [9:0] Pix_604, // sfix10_En0 
 input [9:0] Pix_605, // sfix10_En0 
 input [9:0] Pix_606, // sfix10_En0 
 input [9:0] Pix_607, // sfix10_En0 
 input [9:0] Pix_608, // sfix10_En0 
 input [9:0] Pix_609, // sfix10_En0 
 input [9:0] Pix_610, // sfix10_En0 
 input [9:0] Pix_611, // sfix10_En0 
 input [9:0] Pix_612, // sfix10_En0 
 input [9:0] Pix_613, // sfix10_En0 
 input [9:0] Pix_614, // sfix10_En0 
 input [9:0] Pix_615, // sfix10_En0 
 input [9:0] Pix_616, // sfix10_En0 
 input [9:0] Pix_617, // sfix10_En0 
 input [9:0] Pix_618, // sfix10_En0 
 input [9:0] Pix_619, // sfix10_En0 
 input [9:0] Pix_620, // sfix10_En0 
 input [9:0] Pix_621, // sfix10_En0 
 input [9:0] Pix_622, // sfix10_En0 
 input [9:0] Pix_623, // sfix10_En0 
 input [9:0] Pix_624, // sfix10_En0 
 input [9:0] Pix_625, // sfix10_En0 
 input [9:0] Pix_626, // sfix10_En0 
 input [9:0] Pix_627, // sfix10_En0 
 input [9:0] Pix_628, // sfix10_En0 
 input [9:0] Pix_629, // sfix10_En0 
 input [9:0] Pix_630, // sfix10_En0 
 input [9:0] Pix_631, // sfix10_En0 
 input [9:0] Pix_632, // sfix10_En0 
 input [9:0] Pix_633, // sfix10_En0 
 input [9:0] Pix_634, // sfix10_En0 
 input [9:0] Pix_635, // sfix10_En0 
 input [9:0] Pix_636, // sfix10_En0 
 input [9:0] Pix_637, // sfix10_En0 
 input [9:0] Pix_638, // sfix10_En0 
 input [9:0] Pix_639, // sfix10_En0 
 input [9:0] Pix_640, // sfix10_En0 
 input [9:0] Pix_641, // sfix10_En0 
 input [9:0] Pix_642, // sfix10_En0 
 input [9:0] Pix_643, // sfix10_En0 
 input [9:0] Pix_644, // sfix10_En0 
 input [9:0] Pix_645, // sfix10_En0 
 input [9:0] Pix_646, // sfix10_En0 
 input [9:0] Pix_647, // sfix10_En0 
 input [9:0] Pix_648, // sfix10_En0 
 input [9:0] Pix_649, // sfix10_En0 
 input [9:0] Pix_650, // sfix10_En0 
 input [9:0] Pix_651, // sfix10_En0 
 input [9:0] Pix_652, // sfix10_En0 
 input [9:0] Pix_653, // sfix10_En0 
 input [9:0] Pix_654, // sfix10_En0 
 input [9:0] Pix_655, // sfix10_En0 
 input [9:0] Pix_656, // sfix10_En0 
 input [9:0] Pix_657, // sfix10_En0 
 input [9:0] Pix_658, // sfix10_En0 
 input [9:0] Pix_659, // sfix10_En0 
 input [9:0] Pix_660, // sfix10_En0 
 input [9:0] Pix_661, // sfix10_En0 
 input [9:0] Pix_662, // sfix10_En0 
 input [9:0] Pix_663, // sfix10_En0 
 input [9:0] Pix_664, // sfix10_En0 
 input [9:0] Pix_665, // sfix10_En0 
 input [9:0] Pix_666, // sfix10_En0 
 input [9:0] Pix_667, // sfix10_En0 
 input [9:0] Pix_668, // sfix10_En0 
 input [9:0] Pix_669, // sfix10_En0 
 input [9:0] Pix_670, // sfix10_En0 
 input [9:0] Pix_671, // sfix10_En0 
 input [9:0] Pix_672, // sfix10_En0 
 input [9:0] Pix_673, // sfix10_En0 
 input [9:0] Pix_674, // sfix10_En0 
 input [9:0] Pix_675, // sfix10_En0 
 input [9:0] Pix_676, // sfix10_En0 
 input [9:0] Pix_677, // sfix10_En0 
 input [9:0] Pix_678, // sfix10_En0 
 input [9:0] Pix_679, // sfix10_En0 
 input [9:0] Pix_680, // sfix10_En0 
 input [9:0] Pix_681, // sfix10_En0 
 input [9:0] Pix_682, // sfix10_En0 
 input [9:0] Pix_683, // sfix10_En0 
 input [9:0] Pix_684, // sfix10_En0 
 input [9:0] Pix_685, // sfix10_En0 
 input [9:0] Pix_686, // sfix10_En0 
 input [9:0] Pix_687, // sfix10_En0 
 input [9:0] Pix_688, // sfix10_En0 
 input [9:0] Pix_689, // sfix10_En0 
 input [9:0] Pix_690, // sfix10_En0 
 input [9:0] Pix_691, // sfix10_En0 
 input [9:0] Pix_692, // sfix10_En0 
 input [9:0] Pix_693, // sfix10_En0 
 input [9:0] Pix_694, // sfix10_En0 
 input [9:0] Pix_695, // sfix10_En0 
 input [9:0] Pix_696, // sfix10_En0 
 input [9:0] Pix_697, // sfix10_En0 
 input [9:0] Pix_698, // sfix10_En0 
 input [9:0] Pix_699, // sfix10_En0 
 input [9:0] Pix_700, // sfix10_En0 
 input [9:0] Pix_701, // sfix10_En0 
 input [9:0] Pix_702, // sfix10_En0 
 input [9:0] Pix_703, // sfix10_En0 
 input [9:0] Pix_704, // sfix10_En0 
 input [9:0] Pix_705, // sfix10_En0 
 input [9:0] Pix_706, // sfix10_En0 
 input [9:0] Pix_707, // sfix10_En0 
 input [9:0] Pix_708, // sfix10_En0 
 input [9:0] Pix_709, // sfix10_En0 
 input [9:0] Pix_710, // sfix10_En0 
 input [9:0] Pix_711, // sfix10_En0 
 input [9:0] Pix_712, // sfix10_En0 
 input [9:0] Pix_713, // sfix10_En0 
 input [9:0] Pix_714, // sfix10_En0 
 input [9:0] Pix_715, // sfix10_En0 
 input [9:0] Pix_716, // sfix10_En0 
 input [9:0] Pix_717, // sfix10_En0 
 input [9:0] Pix_718, // sfix10_En0 
 input [9:0] Pix_719, // sfix10_En0 
 input [9:0] Pix_720, // sfix10_En0 
 input [9:0] Pix_721, // sfix10_En0 
 input [9:0] Pix_722, // sfix10_En0 
 input [9:0] Pix_723, // sfix10_En0 
 input [9:0] Pix_724, // sfix10_En0 
 input [9:0] Pix_725, // sfix10_En0 
 input [9:0] Pix_726, // sfix10_En0 
 input [9:0] Pix_727, // sfix10_En0 
 input [9:0] Pix_728, // sfix10_En0 
 input [9:0] Pix_729, // sfix10_En0 
 input [9:0] Pix_730, // sfix10_En0 
 input [9:0] Pix_731, // sfix10_En0 
 input [9:0] Pix_732, // sfix10_En0 
 input [9:0] Pix_733, // sfix10_En0 
 input [9:0] Pix_734, // sfix10_En0 
 input [9:0] Pix_735, // sfix10_En0 
 input [9:0] Pix_736, // sfix10_En0 
 input [9:0] Pix_737, // sfix10_En0 
 input [9:0] Pix_738, // sfix10_En0 
 input [9:0] Pix_739, // sfix10_En0 
 input [9:0] Pix_740, // sfix10_En0 
 input [9:0] Pix_741, // sfix10_En0 
 input [9:0] Pix_742, // sfix10_En0 
 input [9:0] Pix_743, // sfix10_En0 
 input [9:0] Pix_744, // sfix10_En0 
 input [9:0] Pix_745, // sfix10_En0 
 input [9:0] Pix_746, // sfix10_En0 
 input [9:0] Pix_747, // sfix10_En0 
 input [9:0] Pix_748, // sfix10_En0 
 input [9:0] Pix_749, // sfix10_En0 
 input [9:0] Pix_750, // sfix10_En0 
 input [9:0] Pix_751, // sfix10_En0 
 input [9:0] Pix_752, // sfix10_En0 
 input [9:0] Pix_753, // sfix10_En0 
 input [9:0] Pix_754, // sfix10_En0 
 input [9:0] Pix_755, // sfix10_En0 
 input [9:0] Pix_756, // sfix10_En0 
 input [9:0] Pix_757, // sfix10_En0 
 input [9:0] Pix_758, // sfix10_En0 
 input [9:0] Pix_759, // sfix10_En0 
 input [9:0] Pix_760, // sfix10_En0 
 input [9:0] Pix_761, // sfix10_En0 
 input [9:0] Pix_762, // sfix10_En0 
 input [9:0] Pix_763, // sfix10_En0 
 input [9:0] Pix_764, // sfix10_En0 
 input [9:0] Pix_765, // sfix10_En0 
 input [9:0] Pix_766, // sfix10_En0 
 input [9:0] Pix_767, // sfix10_En0 
 input [9:0] Pix_768, // sfix10_En0 
 input [9:0] Pix_769, // sfix10_En0 
 input [9:0] Pix_770, // sfix10_En0 
 input [9:0] Pix_771, // sfix10_En0 
 input [9:0] Pix_772, // sfix10_En0 
 input [9:0] Pix_773, // sfix10_En0 
 input [9:0] Pix_774, // sfix10_En0 
 input [9:0] Pix_775, // sfix10_En0 
 input [9:0] Pix_776, // sfix10_En0 
 input [9:0] Pix_777, // sfix10_En0 
 input [9:0] Pix_778, // sfix10_En0 
 input [9:0] Pix_779, // sfix10_En0 
 input [9:0] Pix_780, // sfix10_En0 
 input [9:0] Pix_781, // sfix10_En0 
 input [9:0] Pix_782, // sfix10_En0 
 input [9:0] Pix_783, // sfix10_En0 
 input [9:0] Pix_784, // sfix10_En0 
 input [18:0] Wgt_0, // sfix19_En18 
  input [18:0] Wgt_1, // sfix19_En18 
  input [18:0] Wgt_2, // sfix19_En18 
  input [18:0] Wgt_3, // sfix19_En18 
  input [18:0] Wgt_4, // sfix19_En18 
  input [18:0] Wgt_5, // sfix19_En18 
  input [18:0] Wgt_6, // sfix19_En18 
  input [18:0] Wgt_7, // sfix19_En18 
  input [18:0] Wgt_8, // sfix19_En18 
  input [18:0] Wgt_9, // sfix19_En18 
  input [18:0] Wgt_10, // sfix19_En18 
  input [18:0] Wgt_11, // sfix19_En18 
  input [18:0] Wgt_12, // sfix19_En18 
  input [18:0] Wgt_13, // sfix19_En18 
  input [18:0] Wgt_14, // sfix19_En18 
  input [18:0] Wgt_15, // sfix19_En18 
  input [18:0] Wgt_16, // sfix19_En18 
  input [18:0] Wgt_17, // sfix19_En18 
  input [18:0] Wgt_18, // sfix19_En18 
  input [18:0] Wgt_19, // sfix19_En18 
  input [18:0] Wgt_20, // sfix19_En18 
  input [18:0] Wgt_21, // sfix19_En18 
  input [18:0] Wgt_22, // sfix19_En18 
  input [18:0] Wgt_23, // sfix19_En18 
  input [18:0] Wgt_24, // sfix19_En18 
  input [18:0] Wgt_25, // sfix19_En18 
  input [18:0] Wgt_26, // sfix19_En18 
  input [18:0] Wgt_27, // sfix19_En18 
  input [18:0] Wgt_28, // sfix19_En18 
  input [18:0] Wgt_29, // sfix19_En18 
  input [18:0] Wgt_30, // sfix19_En18 
  input [18:0] Wgt_31, // sfix19_En18 
  input [18:0] Wgt_32, // sfix19_En18 
  input [18:0] Wgt_33, // sfix19_En18 
  input [18:0] Wgt_34, // sfix19_En18 
  input [18:0] Wgt_35, // sfix19_En18 
  input [18:0] Wgt_36, // sfix19_En18 
  input [18:0] Wgt_37, // sfix19_En18 
  input [18:0] Wgt_38, // sfix19_En18 
  input [18:0] Wgt_39, // sfix19_En18 
  input [18:0] Wgt_40, // sfix19_En18 
  input [18:0] Wgt_41, // sfix19_En18 
  input [18:0] Wgt_42, // sfix19_En18 
  input [18:0] Wgt_43, // sfix19_En18 
  input [18:0] Wgt_44, // sfix19_En18 
  input [18:0] Wgt_45, // sfix19_En18 
  input [18:0] Wgt_46, // sfix19_En18 
  input [18:0] Wgt_47, // sfix19_En18 
  input [18:0] Wgt_48, // sfix19_En18 
  input [18:0] Wgt_49, // sfix19_En18 
  input [18:0] Wgt_50, // sfix19_En18 
  input [18:0] Wgt_51, // sfix19_En18 
  input [18:0] Wgt_52, // sfix19_En18 
  input [18:0] Wgt_53, // sfix19_En18 
  input [18:0] Wgt_54, // sfix19_En18 
  input [18:0] Wgt_55, // sfix19_En18 
  input [18:0] Wgt_56, // sfix19_En18 
  input [18:0] Wgt_57, // sfix19_En18 
  input [18:0] Wgt_58, // sfix19_En18 
  input [18:0] Wgt_59, // sfix19_En18 
  input [18:0] Wgt_60, // sfix19_En18 
  input [18:0] Wgt_61, // sfix19_En18 
  input [18:0] Wgt_62, // sfix19_En18 
  input [18:0] Wgt_63, // sfix19_En18 
  input [18:0] Wgt_64, // sfix19_En18 
  input [18:0] Wgt_65, // sfix19_En18 
  input [18:0] Wgt_66, // sfix19_En18 
  input [18:0] Wgt_67, // sfix19_En18 
  input [18:0] Wgt_68, // sfix19_En18 
  input [18:0] Wgt_69, // sfix19_En18 
  input [18:0] Wgt_70, // sfix19_En18 
  input [18:0] Wgt_71, // sfix19_En18 
  input [18:0] Wgt_72, // sfix19_En18 
  input [18:0] Wgt_73, // sfix19_En18 
  input [18:0] Wgt_74, // sfix19_En18 
  input [18:0] Wgt_75, // sfix19_En18 
  input [18:0] Wgt_76, // sfix19_En18 
  input [18:0] Wgt_77, // sfix19_En18 
  input [18:0] Wgt_78, // sfix19_En18 
  input [18:0] Wgt_79, // sfix19_En18 
  input [18:0] Wgt_80, // sfix19_En18 
  input [18:0] Wgt_81, // sfix19_En18 
  input [18:0] Wgt_82, // sfix19_En18 
  input [18:0] Wgt_83, // sfix19_En18 
  input [18:0] Wgt_84, // sfix19_En18 
  input [18:0] Wgt_85, // sfix19_En18 
  input [18:0] Wgt_86, // sfix19_En18 
  input [18:0] Wgt_87, // sfix19_En18 
  input [18:0] Wgt_88, // sfix19_En18 
  input [18:0] Wgt_89, // sfix19_En18 
  input [18:0] Wgt_90, // sfix19_En18 
  input [18:0] Wgt_91, // sfix19_En18 
  input [18:0] Wgt_92, // sfix19_En18 
  input [18:0] Wgt_93, // sfix19_En18 
  input [18:0] Wgt_94, // sfix19_En18 
  input [18:0] Wgt_95, // sfix19_En18 
  input [18:0] Wgt_96, // sfix19_En18 
  input [18:0] Wgt_97, // sfix19_En18 
  input [18:0] Wgt_98, // sfix19_En18 
  input [18:0] Wgt_99, // sfix19_En18 
  input [18:0] Wgt_100, // sfix19_En18 
  input [18:0] Wgt_101, // sfix19_En18 
  input [18:0] Wgt_102, // sfix19_En18 
  input [18:0] Wgt_103, // sfix19_En18 
  input [18:0] Wgt_104, // sfix19_En18 
  input [18:0] Wgt_105, // sfix19_En18 
  input [18:0] Wgt_106, // sfix19_En18 
  input [18:0] Wgt_107, // sfix19_En18 
  input [18:0] Wgt_108, // sfix19_En18 
  input [18:0] Wgt_109, // sfix19_En18 
  input [18:0] Wgt_110, // sfix19_En18 
  input [18:0] Wgt_111, // sfix19_En18 
  input [18:0] Wgt_112, // sfix19_En18 
  input [18:0] Wgt_113, // sfix19_En18 
  input [18:0] Wgt_114, // sfix19_En18 
  input [18:0] Wgt_115, // sfix19_En18 
  input [18:0] Wgt_116, // sfix19_En18 
  input [18:0] Wgt_117, // sfix19_En18 
  input [18:0] Wgt_118, // sfix19_En18 
  input [18:0] Wgt_119, // sfix19_En18 
  input [18:0] Wgt_120, // sfix19_En18 
  input [18:0] Wgt_121, // sfix19_En18 
  input [18:0] Wgt_122, // sfix19_En18 
  input [18:0] Wgt_123, // sfix19_En18 
  input [18:0] Wgt_124, // sfix19_En18 
  input [18:0] Wgt_125, // sfix19_En18 
  input [18:0] Wgt_126, // sfix19_En18 
  input [18:0] Wgt_127, // sfix19_En18 
  input [18:0] Wgt_128, // sfix19_En18 
  input [18:0] Wgt_129, // sfix19_En18 
  input [18:0] Wgt_130, // sfix19_En18 
  input [18:0] Wgt_131, // sfix19_En18 
  input [18:0] Wgt_132, // sfix19_En18 
  input [18:0] Wgt_133, // sfix19_En18 
  input [18:0] Wgt_134, // sfix19_En18 
  input [18:0] Wgt_135, // sfix19_En18 
  input [18:0] Wgt_136, // sfix19_En18 
  input [18:0] Wgt_137, // sfix19_En18 
  input [18:0] Wgt_138, // sfix19_En18 
  input [18:0] Wgt_139, // sfix19_En18 
  input [18:0] Wgt_140, // sfix19_En18 
  input [18:0] Wgt_141, // sfix19_En18 
  input [18:0] Wgt_142, // sfix19_En18 
  input [18:0] Wgt_143, // sfix19_En18 
  input [18:0] Wgt_144, // sfix19_En18 
  input [18:0] Wgt_145, // sfix19_En18 
  input [18:0] Wgt_146, // sfix19_En18 
  input [18:0] Wgt_147, // sfix19_En18 
  input [18:0] Wgt_148, // sfix19_En18 
  input [18:0] Wgt_149, // sfix19_En18 
  input [18:0] Wgt_150, // sfix19_En18 
  input [18:0] Wgt_151, // sfix19_En18 
  input [18:0] Wgt_152, // sfix19_En18 
  input [18:0] Wgt_153, // sfix19_En18 
  input [18:0] Wgt_154, // sfix19_En18 
  input [18:0] Wgt_155, // sfix19_En18 
  input [18:0] Wgt_156, // sfix19_En18 
  input [18:0] Wgt_157, // sfix19_En18 
  input [18:0] Wgt_158, // sfix19_En18 
  input [18:0] Wgt_159, // sfix19_En18 
  input [18:0] Wgt_160, // sfix19_En18 
  input [18:0] Wgt_161, // sfix19_En18 
  input [18:0] Wgt_162, // sfix19_En18 
  input [18:0] Wgt_163, // sfix19_En18 
  input [18:0] Wgt_164, // sfix19_En18 
  input [18:0] Wgt_165, // sfix19_En18 
  input [18:0] Wgt_166, // sfix19_En18 
  input [18:0] Wgt_167, // sfix19_En18 
  input [18:0] Wgt_168, // sfix19_En18 
  input [18:0] Wgt_169, // sfix19_En18 
  input [18:0] Wgt_170, // sfix19_En18 
  input [18:0] Wgt_171, // sfix19_En18 
  input [18:0] Wgt_172, // sfix19_En18 
  input [18:0] Wgt_173, // sfix19_En18 
  input [18:0] Wgt_174, // sfix19_En18 
  input [18:0] Wgt_175, // sfix19_En18 
  input [18:0] Wgt_176, // sfix19_En18 
  input [18:0] Wgt_177, // sfix19_En18 
  input [18:0] Wgt_178, // sfix19_En18 
  input [18:0] Wgt_179, // sfix19_En18 
  input [18:0] Wgt_180, // sfix19_En18 
  input [18:0] Wgt_181, // sfix19_En18 
  input [18:0] Wgt_182, // sfix19_En18 
  input [18:0] Wgt_183, // sfix19_En18 
  input [18:0] Wgt_184, // sfix19_En18 
  input [18:0] Wgt_185, // sfix19_En18 
  input [18:0] Wgt_186, // sfix19_En18 
  input [18:0] Wgt_187, // sfix19_En18 
  input [18:0] Wgt_188, // sfix19_En18 
  input [18:0] Wgt_189, // sfix19_En18 
  input [18:0] Wgt_190, // sfix19_En18 
  input [18:0] Wgt_191, // sfix19_En18 
  input [18:0] Wgt_192, // sfix19_En18 
  input [18:0] Wgt_193, // sfix19_En18 
  input [18:0] Wgt_194, // sfix19_En18 
  input [18:0] Wgt_195, // sfix19_En18 
  input [18:0] Wgt_196, // sfix19_En18 
  input [18:0] Wgt_197, // sfix19_En18 
  input [18:0] Wgt_198, // sfix19_En18 
  input [18:0] Wgt_199, // sfix19_En18 
  input [18:0] Wgt_200, // sfix19_En18 
  input [18:0] Wgt_201, // sfix19_En18 
  input [18:0] Wgt_202, // sfix19_En18 
  input [18:0] Wgt_203, // sfix19_En18 
  input [18:0] Wgt_204, // sfix19_En18 
  input [18:0] Wgt_205, // sfix19_En18 
  input [18:0] Wgt_206, // sfix19_En18 
  input [18:0] Wgt_207, // sfix19_En18 
  input [18:0] Wgt_208, // sfix19_En18 
  input [18:0] Wgt_209, // sfix19_En18 
  input [18:0] Wgt_210, // sfix19_En18 
  input [18:0] Wgt_211, // sfix19_En18 
  input [18:0] Wgt_212, // sfix19_En18 
  input [18:0] Wgt_213, // sfix19_En18 
  input [18:0] Wgt_214, // sfix19_En18 
  input [18:0] Wgt_215, // sfix19_En18 
  input [18:0] Wgt_216, // sfix19_En18 
  input [18:0] Wgt_217, // sfix19_En18 
  input [18:0] Wgt_218, // sfix19_En18 
  input [18:0] Wgt_219, // sfix19_En18 
  input [18:0] Wgt_220, // sfix19_En18 
  input [18:0] Wgt_221, // sfix19_En18 
  input [18:0] Wgt_222, // sfix19_En18 
  input [18:0] Wgt_223, // sfix19_En18 
  input [18:0] Wgt_224, // sfix19_En18 
  input [18:0] Wgt_225, // sfix19_En18 
  input [18:0] Wgt_226, // sfix19_En18 
  input [18:0] Wgt_227, // sfix19_En18 
  input [18:0] Wgt_228, // sfix19_En18 
  input [18:0] Wgt_229, // sfix19_En18 
  input [18:0] Wgt_230, // sfix19_En18 
  input [18:0] Wgt_231, // sfix19_En18 
  input [18:0] Wgt_232, // sfix19_En18 
  input [18:0] Wgt_233, // sfix19_En18 
  input [18:0] Wgt_234, // sfix19_En18 
  input [18:0] Wgt_235, // sfix19_En18 
  input [18:0] Wgt_236, // sfix19_En18 
  input [18:0] Wgt_237, // sfix19_En18 
  input [18:0] Wgt_238, // sfix19_En18 
  input [18:0] Wgt_239, // sfix19_En18 
  input [18:0] Wgt_240, // sfix19_En18 
  input [18:0] Wgt_241, // sfix19_En18 
  input [18:0] Wgt_242, // sfix19_En18 
  input [18:0] Wgt_243, // sfix19_En18 
  input [18:0] Wgt_244, // sfix19_En18 
  input [18:0] Wgt_245, // sfix19_En18 
  input [18:0] Wgt_246, // sfix19_En18 
  input [18:0] Wgt_247, // sfix19_En18 
  input [18:0] Wgt_248, // sfix19_En18 
  input [18:0] Wgt_249, // sfix19_En18 
  input [18:0] Wgt_250, // sfix19_En18 
  input [18:0] Wgt_251, // sfix19_En18 
  input [18:0] Wgt_252, // sfix19_En18 
  input [18:0] Wgt_253, // sfix19_En18 
  input [18:0] Wgt_254, // sfix19_En18 
  input [18:0] Wgt_255, // sfix19_En18 
  input [18:0] Wgt_256, // sfix19_En18 
  input [18:0] Wgt_257, // sfix19_En18 
  input [18:0] Wgt_258, // sfix19_En18 
  input [18:0] Wgt_259, // sfix19_En18 
  input [18:0] Wgt_260, // sfix19_En18 
  input [18:0] Wgt_261, // sfix19_En18 
  input [18:0] Wgt_262, // sfix19_En18 
  input [18:0] Wgt_263, // sfix19_En18 
  input [18:0] Wgt_264, // sfix19_En18 
  input [18:0] Wgt_265, // sfix19_En18 
  input [18:0] Wgt_266, // sfix19_En18 
  input [18:0] Wgt_267, // sfix19_En18 
  input [18:0] Wgt_268, // sfix19_En18 
  input [18:0] Wgt_269, // sfix19_En18 
  input [18:0] Wgt_270, // sfix19_En18 
  input [18:0] Wgt_271, // sfix19_En18 
  input [18:0] Wgt_272, // sfix19_En18 
  input [18:0] Wgt_273, // sfix19_En18 
  input [18:0] Wgt_274, // sfix19_En18 
  input [18:0] Wgt_275, // sfix19_En18 
  input [18:0] Wgt_276, // sfix19_En18 
  input [18:0] Wgt_277, // sfix19_En18 
  input [18:0] Wgt_278, // sfix19_En18 
  input [18:0] Wgt_279, // sfix19_En18 
  input [18:0] Wgt_280, // sfix19_En18 
  input [18:0] Wgt_281, // sfix19_En18 
  input [18:0] Wgt_282, // sfix19_En18 
  input [18:0] Wgt_283, // sfix19_En18 
  input [18:0] Wgt_284, // sfix19_En18 
  input [18:0] Wgt_285, // sfix19_En18 
  input [18:0] Wgt_286, // sfix19_En18 
  input [18:0] Wgt_287, // sfix19_En18 
  input [18:0] Wgt_288, // sfix19_En18 
  input [18:0] Wgt_289, // sfix19_En18 
  input [18:0] Wgt_290, // sfix19_En18 
  input [18:0] Wgt_291, // sfix19_En18 
  input [18:0] Wgt_292, // sfix19_En18 
  input [18:0] Wgt_293, // sfix19_En18 
  input [18:0] Wgt_294, // sfix19_En18 
  input [18:0] Wgt_295, // sfix19_En18 
  input [18:0] Wgt_296, // sfix19_En18 
  input [18:0] Wgt_297, // sfix19_En18 
  input [18:0] Wgt_298, // sfix19_En18 
  input [18:0] Wgt_299, // sfix19_En18 
  input [18:0] Wgt_300, // sfix19_En18 
  input [18:0] Wgt_301, // sfix19_En18 
  input [18:0] Wgt_302, // sfix19_En18 
  input [18:0] Wgt_303, // sfix19_En18 
  input [18:0] Wgt_304, // sfix19_En18 
  input [18:0] Wgt_305, // sfix19_En18 
  input [18:0] Wgt_306, // sfix19_En18 
  input [18:0] Wgt_307, // sfix19_En18 
  input [18:0] Wgt_308, // sfix19_En18 
  input [18:0] Wgt_309, // sfix19_En18 
  input [18:0] Wgt_310, // sfix19_En18 
  input [18:0] Wgt_311, // sfix19_En18 
  input [18:0] Wgt_312, // sfix19_En18 
  input [18:0] Wgt_313, // sfix19_En18 
  input [18:0] Wgt_314, // sfix19_En18 
  input [18:0] Wgt_315, // sfix19_En18 
  input [18:0] Wgt_316, // sfix19_En18 
  input [18:0] Wgt_317, // sfix19_En18 
  input [18:0] Wgt_318, // sfix19_En18 
  input [18:0] Wgt_319, // sfix19_En18 
  input [18:0] Wgt_320, // sfix19_En18 
  input [18:0] Wgt_321, // sfix19_En18 
  input [18:0] Wgt_322, // sfix19_En18 
  input [18:0] Wgt_323, // sfix19_En18 
  input [18:0] Wgt_324, // sfix19_En18 
  input [18:0] Wgt_325, // sfix19_En18 
  input [18:0] Wgt_326, // sfix19_En18 
  input [18:0] Wgt_327, // sfix19_En18 
  input [18:0] Wgt_328, // sfix19_En18 
  input [18:0] Wgt_329, // sfix19_En18 
  input [18:0] Wgt_330, // sfix19_En18 
  input [18:0] Wgt_331, // sfix19_En18 
  input [18:0] Wgt_332, // sfix19_En18 
  input [18:0] Wgt_333, // sfix19_En18 
  input [18:0] Wgt_334, // sfix19_En18 
  input [18:0] Wgt_335, // sfix19_En18 
  input [18:0] Wgt_336, // sfix19_En18 
  input [18:0] Wgt_337, // sfix19_En18 
  input [18:0] Wgt_338, // sfix19_En18 
  input [18:0] Wgt_339, // sfix19_En18 
  input [18:0] Wgt_340, // sfix19_En18 
  input [18:0] Wgt_341, // sfix19_En18 
  input [18:0] Wgt_342, // sfix19_En18 
  input [18:0] Wgt_343, // sfix19_En18 
  input [18:0] Wgt_344, // sfix19_En18 
  input [18:0] Wgt_345, // sfix19_En18 
  input [18:0] Wgt_346, // sfix19_En18 
  input [18:0] Wgt_347, // sfix19_En18 
  input [18:0] Wgt_348, // sfix19_En18 
  input [18:0] Wgt_349, // sfix19_En18 
  input [18:0] Wgt_350, // sfix19_En18 
  input [18:0] Wgt_351, // sfix19_En18 
  input [18:0] Wgt_352, // sfix19_En18 
  input [18:0] Wgt_353, // sfix19_En18 
  input [18:0] Wgt_354, // sfix19_En18 
  input [18:0] Wgt_355, // sfix19_En18 
  input [18:0] Wgt_356, // sfix19_En18 
  input [18:0] Wgt_357, // sfix19_En18 
  input [18:0] Wgt_358, // sfix19_En18 
  input [18:0] Wgt_359, // sfix19_En18 
  input [18:0] Wgt_360, // sfix19_En18 
  input [18:0] Wgt_361, // sfix19_En18 
  input [18:0] Wgt_362, // sfix19_En18 
  input [18:0] Wgt_363, // sfix19_En18 
  input [18:0] Wgt_364, // sfix19_En18 
  input [18:0] Wgt_365, // sfix19_En18 
  input [18:0] Wgt_366, // sfix19_En18 
  input [18:0] Wgt_367, // sfix19_En18 
  input [18:0] Wgt_368, // sfix19_En18 
  input [18:0] Wgt_369, // sfix19_En18 
  input [18:0] Wgt_370, // sfix19_En18 
  input [18:0] Wgt_371, // sfix19_En18 
  input [18:0] Wgt_372, // sfix19_En18 
  input [18:0] Wgt_373, // sfix19_En18 
  input [18:0] Wgt_374, // sfix19_En18 
  input [18:0] Wgt_375, // sfix19_En18 
  input [18:0] Wgt_376, // sfix19_En18 
  input [18:0] Wgt_377, // sfix19_En18 
  input [18:0] Wgt_378, // sfix19_En18 
  input [18:0] Wgt_379, // sfix19_En18 
  input [18:0] Wgt_380, // sfix19_En18 
  input [18:0] Wgt_381, // sfix19_En18 
  input [18:0] Wgt_382, // sfix19_En18 
  input [18:0] Wgt_383, // sfix19_En18 
  input [18:0] Wgt_384, // sfix19_En18 
  input [18:0] Wgt_385, // sfix19_En18 
  input [18:0] Wgt_386, // sfix19_En18 
  input [18:0] Wgt_387, // sfix19_En18 
  input [18:0] Wgt_388, // sfix19_En18 
  input [18:0] Wgt_389, // sfix19_En18 
  input [18:0] Wgt_390, // sfix19_En18 
  input [18:0] Wgt_391, // sfix19_En18 
  input [18:0] Wgt_392, // sfix19_En18 
  input [18:0] Wgt_393, // sfix19_En18 
  input [18:0] Wgt_394, // sfix19_En18 
  input [18:0] Wgt_395, // sfix19_En18 
  input [18:0] Wgt_396, // sfix19_En18 
  input [18:0] Wgt_397, // sfix19_En18 
  input [18:0] Wgt_398, // sfix19_En18 
  input [18:0] Wgt_399, // sfix19_En18 
  input [18:0] Wgt_400, // sfix19_En18 
  input [18:0] Wgt_401, // sfix19_En18 
  input [18:0] Wgt_402, // sfix19_En18 
  input [18:0] Wgt_403, // sfix19_En18 
  input [18:0] Wgt_404, // sfix19_En18 
  input [18:0] Wgt_405, // sfix19_En18 
  input [18:0] Wgt_406, // sfix19_En18 
  input [18:0] Wgt_407, // sfix19_En18 
  input [18:0] Wgt_408, // sfix19_En18 
  input [18:0] Wgt_409, // sfix19_En18 
  input [18:0] Wgt_410, // sfix19_En18 
  input [18:0] Wgt_411, // sfix19_En18 
  input [18:0] Wgt_412, // sfix19_En18 
  input [18:0] Wgt_413, // sfix19_En18 
  input [18:0] Wgt_414, // sfix19_En18 
  input [18:0] Wgt_415, // sfix19_En18 
  input [18:0] Wgt_416, // sfix19_En18 
  input [18:0] Wgt_417, // sfix19_En18 
  input [18:0] Wgt_418, // sfix19_En18 
  input [18:0] Wgt_419, // sfix19_En18 
  input [18:0] Wgt_420, // sfix19_En18 
  input [18:0] Wgt_421, // sfix19_En18 
  input [18:0] Wgt_422, // sfix19_En18 
  input [18:0] Wgt_423, // sfix19_En18 
  input [18:0] Wgt_424, // sfix19_En18 
  input [18:0] Wgt_425, // sfix19_En18 
  input [18:0] Wgt_426, // sfix19_En18 
  input [18:0] Wgt_427, // sfix19_En18 
  input [18:0] Wgt_428, // sfix19_En18 
  input [18:0] Wgt_429, // sfix19_En18 
  input [18:0] Wgt_430, // sfix19_En18 
  input [18:0] Wgt_431, // sfix19_En18 
  input [18:0] Wgt_432, // sfix19_En18 
  input [18:0] Wgt_433, // sfix19_En18 
  input [18:0] Wgt_434, // sfix19_En18 
  input [18:0] Wgt_435, // sfix19_En18 
  input [18:0] Wgt_436, // sfix19_En18 
  input [18:0] Wgt_437, // sfix19_En18 
  input [18:0] Wgt_438, // sfix19_En18 
  input [18:0] Wgt_439, // sfix19_En18 
  input [18:0] Wgt_440, // sfix19_En18 
  input [18:0] Wgt_441, // sfix19_En18 
  input [18:0] Wgt_442, // sfix19_En18 
  input [18:0] Wgt_443, // sfix19_En18 
  input [18:0] Wgt_444, // sfix19_En18 
  input [18:0] Wgt_445, // sfix19_En18 
  input [18:0] Wgt_446, // sfix19_En18 
  input [18:0] Wgt_447, // sfix19_En18 
  input [18:0] Wgt_448, // sfix19_En18 
  input [18:0] Wgt_449, // sfix19_En18 
  input [18:0] Wgt_450, // sfix19_En18 
  input [18:0] Wgt_451, // sfix19_En18 
  input [18:0] Wgt_452, // sfix19_En18 
  input [18:0] Wgt_453, // sfix19_En18 
  input [18:0] Wgt_454, // sfix19_En18 
  input [18:0] Wgt_455, // sfix19_En18 
  input [18:0] Wgt_456, // sfix19_En18 
  input [18:0] Wgt_457, // sfix19_En18 
  input [18:0] Wgt_458, // sfix19_En18 
  input [18:0] Wgt_459, // sfix19_En18 
  input [18:0] Wgt_460, // sfix19_En18 
  input [18:0] Wgt_461, // sfix19_En18 
  input [18:0] Wgt_462, // sfix19_En18 
  input [18:0] Wgt_463, // sfix19_En18 
  input [18:0] Wgt_464, // sfix19_En18 
  input [18:0] Wgt_465, // sfix19_En18 
  input [18:0] Wgt_466, // sfix19_En18 
  input [18:0] Wgt_467, // sfix19_En18 
  input [18:0] Wgt_468, // sfix19_En18 
  input [18:0] Wgt_469, // sfix19_En18 
  input [18:0] Wgt_470, // sfix19_En18 
  input [18:0] Wgt_471, // sfix19_En18 
  input [18:0] Wgt_472, // sfix19_En18 
  input [18:0] Wgt_473, // sfix19_En18 
  input [18:0] Wgt_474, // sfix19_En18 
  input [18:0] Wgt_475, // sfix19_En18 
  input [18:0] Wgt_476, // sfix19_En18 
  input [18:0] Wgt_477, // sfix19_En18 
  input [18:0] Wgt_478, // sfix19_En18 
  input [18:0] Wgt_479, // sfix19_En18 
  input [18:0] Wgt_480, // sfix19_En18 
  input [18:0] Wgt_481, // sfix19_En18 
  input [18:0] Wgt_482, // sfix19_En18 
  input [18:0] Wgt_483, // sfix19_En18 
  input [18:0] Wgt_484, // sfix19_En18 
  input [18:0] Wgt_485, // sfix19_En18 
  input [18:0] Wgt_486, // sfix19_En18 
  input [18:0] Wgt_487, // sfix19_En18 
  input [18:0] Wgt_488, // sfix19_En18 
  input [18:0] Wgt_489, // sfix19_En18 
  input [18:0] Wgt_490, // sfix19_En18 
  input [18:0] Wgt_491, // sfix19_En18 
  input [18:0] Wgt_492, // sfix19_En18 
  input [18:0] Wgt_493, // sfix19_En18 
  input [18:0] Wgt_494, // sfix19_En18 
  input [18:0] Wgt_495, // sfix19_En18 
  input [18:0] Wgt_496, // sfix19_En18 
  input [18:0] Wgt_497, // sfix19_En18 
  input [18:0] Wgt_498, // sfix19_En18 
  input [18:0] Wgt_499, // sfix19_En18 
  input [18:0] Wgt_500, // sfix19_En18 
  input [18:0] Wgt_501, // sfix19_En18 
  input [18:0] Wgt_502, // sfix19_En18 
  input [18:0] Wgt_503, // sfix19_En18 
  input [18:0] Wgt_504, // sfix19_En18 
  input [18:0] Wgt_505, // sfix19_En18 
  input [18:0] Wgt_506, // sfix19_En18 
  input [18:0] Wgt_507, // sfix19_En18 
  input [18:0] Wgt_508, // sfix19_En18 
  input [18:0] Wgt_509, // sfix19_En18 
  input [18:0] Wgt_510, // sfix19_En18 
  input [18:0] Wgt_511, // sfix19_En18 
  input [18:0] Wgt_512, // sfix19_En18 
  input [18:0] Wgt_513, // sfix19_En18 
  input [18:0] Wgt_514, // sfix19_En18 
  input [18:0] Wgt_515, // sfix19_En18 
  input [18:0] Wgt_516, // sfix19_En18 
  input [18:0] Wgt_517, // sfix19_En18 
  input [18:0] Wgt_518, // sfix19_En18 
  input [18:0] Wgt_519, // sfix19_En18 
  input [18:0] Wgt_520, // sfix19_En18 
  input [18:0] Wgt_521, // sfix19_En18 
  input [18:0] Wgt_522, // sfix19_En18 
  input [18:0] Wgt_523, // sfix19_En18 
  input [18:0] Wgt_524, // sfix19_En18 
  input [18:0] Wgt_525, // sfix19_En18 
  input [18:0] Wgt_526, // sfix19_En18 
  input [18:0] Wgt_527, // sfix19_En18 
  input [18:0] Wgt_528, // sfix19_En18 
  input [18:0] Wgt_529, // sfix19_En18 
  input [18:0] Wgt_530, // sfix19_En18 
  input [18:0] Wgt_531, // sfix19_En18 
  input [18:0] Wgt_532, // sfix19_En18 
  input [18:0] Wgt_533, // sfix19_En18 
  input [18:0] Wgt_534, // sfix19_En18 
  input [18:0] Wgt_535, // sfix19_En18 
  input [18:0] Wgt_536, // sfix19_En18 
  input [18:0] Wgt_537, // sfix19_En18 
  input [18:0] Wgt_538, // sfix19_En18 
  input [18:0] Wgt_539, // sfix19_En18 
  input [18:0] Wgt_540, // sfix19_En18 
  input [18:0] Wgt_541, // sfix19_En18 
  input [18:0] Wgt_542, // sfix19_En18 
  input [18:0] Wgt_543, // sfix19_En18 
  input [18:0] Wgt_544, // sfix19_En18 
  input [18:0] Wgt_545, // sfix19_En18 
  input [18:0] Wgt_546, // sfix19_En18 
  input [18:0] Wgt_547, // sfix19_En18 
  input [18:0] Wgt_548, // sfix19_En18 
  input [18:0] Wgt_549, // sfix19_En18 
  input [18:0] Wgt_550, // sfix19_En18 
  input [18:0] Wgt_551, // sfix19_En18 
  input [18:0] Wgt_552, // sfix19_En18 
  input [18:0] Wgt_553, // sfix19_En18 
  input [18:0] Wgt_554, // sfix19_En18 
  input [18:0] Wgt_555, // sfix19_En18 
  input [18:0] Wgt_556, // sfix19_En18 
  input [18:0] Wgt_557, // sfix19_En18 
  input [18:0] Wgt_558, // sfix19_En18 
  input [18:0] Wgt_559, // sfix19_En18 
  input [18:0] Wgt_560, // sfix19_En18 
  input [18:0] Wgt_561, // sfix19_En18 
  input [18:0] Wgt_562, // sfix19_En18 
  input [18:0] Wgt_563, // sfix19_En18 
  input [18:0] Wgt_564, // sfix19_En18 
  input [18:0] Wgt_565, // sfix19_En18 
  input [18:0] Wgt_566, // sfix19_En18 
  input [18:0] Wgt_567, // sfix19_En18 
  input [18:0] Wgt_568, // sfix19_En18 
  input [18:0] Wgt_569, // sfix19_En18 
  input [18:0] Wgt_570, // sfix19_En18 
  input [18:0] Wgt_571, // sfix19_En18 
  input [18:0] Wgt_572, // sfix19_En18 
  input [18:0] Wgt_573, // sfix19_En18 
  input [18:0] Wgt_574, // sfix19_En18 
  input [18:0] Wgt_575, // sfix19_En18 
  input [18:0] Wgt_576, // sfix19_En18 
  input [18:0] Wgt_577, // sfix19_En18 
  input [18:0] Wgt_578, // sfix19_En18 
  input [18:0] Wgt_579, // sfix19_En18 
  input [18:0] Wgt_580, // sfix19_En18 
  input [18:0] Wgt_581, // sfix19_En18 
  input [18:0] Wgt_582, // sfix19_En18 
  input [18:0] Wgt_583, // sfix19_En18 
  input [18:0] Wgt_584, // sfix19_En18 
  input [18:0] Wgt_585, // sfix19_En18 
  input [18:0] Wgt_586, // sfix19_En18 
  input [18:0] Wgt_587, // sfix19_En18 
  input [18:0] Wgt_588, // sfix19_En18 
  input [18:0] Wgt_589, // sfix19_En18 
  input [18:0] Wgt_590, // sfix19_En18 
  input [18:0] Wgt_591, // sfix19_En18 
  input [18:0] Wgt_592, // sfix19_En18 
  input [18:0] Wgt_593, // sfix19_En18 
  input [18:0] Wgt_594, // sfix19_En18 
  input [18:0] Wgt_595, // sfix19_En18 
  input [18:0] Wgt_596, // sfix19_En18 
  input [18:0] Wgt_597, // sfix19_En18 
  input [18:0] Wgt_598, // sfix19_En18 
  input [18:0] Wgt_599, // sfix19_En18 
  input [18:0] Wgt_600, // sfix19_En18 
  input [18:0] Wgt_601, // sfix19_En18 
  input [18:0] Wgt_602, // sfix19_En18 
  input [18:0] Wgt_603, // sfix19_En18 
  input [18:0] Wgt_604, // sfix19_En18 
  input [18:0] Wgt_605, // sfix19_En18 
  input [18:0] Wgt_606, // sfix19_En18 
  input [18:0] Wgt_607, // sfix19_En18 
  input [18:0] Wgt_608, // sfix19_En18 
  input [18:0] Wgt_609, // sfix19_En18 
  input [18:0] Wgt_610, // sfix19_En18 
  input [18:0] Wgt_611, // sfix19_En18 
  input [18:0] Wgt_612, // sfix19_En18 
  input [18:0] Wgt_613, // sfix19_En18 
  input [18:0] Wgt_614, // sfix19_En18 
  input [18:0] Wgt_615, // sfix19_En18 
  input [18:0] Wgt_616, // sfix19_En18 
  input [18:0] Wgt_617, // sfix19_En18 
  input [18:0] Wgt_618, // sfix19_En18 
  input [18:0] Wgt_619, // sfix19_En18 
  input [18:0] Wgt_620, // sfix19_En18 
  input [18:0] Wgt_621, // sfix19_En18 
  input [18:0] Wgt_622, // sfix19_En18 
  input [18:0] Wgt_623, // sfix19_En18 
  input [18:0] Wgt_624, // sfix19_En18 
  input [18:0] Wgt_625, // sfix19_En18 
  input [18:0] Wgt_626, // sfix19_En18 
  input [18:0] Wgt_627, // sfix19_En18 
  input [18:0] Wgt_628, // sfix19_En18 
  input [18:0] Wgt_629, // sfix19_En18 
  input [18:0] Wgt_630, // sfix19_En18 
  input [18:0] Wgt_631, // sfix19_En18 
  input [18:0] Wgt_632, // sfix19_En18 
  input [18:0] Wgt_633, // sfix19_En18 
  input [18:0] Wgt_634, // sfix19_En18 
  input [18:0] Wgt_635, // sfix19_En18 
  input [18:0] Wgt_636, // sfix19_En18 
  input [18:0] Wgt_637, // sfix19_En18 
  input [18:0] Wgt_638, // sfix19_En18 
  input [18:0] Wgt_639, // sfix19_En18 
  input [18:0] Wgt_640, // sfix19_En18 
  input [18:0] Wgt_641, // sfix19_En18 
  input [18:0] Wgt_642, // sfix19_En18 
  input [18:0] Wgt_643, // sfix19_En18 
  input [18:0] Wgt_644, // sfix19_En18 
  input [18:0] Wgt_645, // sfix19_En18 
  input [18:0] Wgt_646, // sfix19_En18 
  input [18:0] Wgt_647, // sfix19_En18 
  input [18:0] Wgt_648, // sfix19_En18 
  input [18:0] Wgt_649, // sfix19_En18 
  input [18:0] Wgt_650, // sfix19_En18 
  input [18:0] Wgt_651, // sfix19_En18 
  input [18:0] Wgt_652, // sfix19_En18 
  input [18:0] Wgt_653, // sfix19_En18 
  input [18:0] Wgt_654, // sfix19_En18 
  input [18:0] Wgt_655, // sfix19_En18 
  input [18:0] Wgt_656, // sfix19_En18 
  input [18:0] Wgt_657, // sfix19_En18 
  input [18:0] Wgt_658, // sfix19_En18 
  input [18:0] Wgt_659, // sfix19_En18 
  input [18:0] Wgt_660, // sfix19_En18 
  input [18:0] Wgt_661, // sfix19_En18 
  input [18:0] Wgt_662, // sfix19_En18 
  input [18:0] Wgt_663, // sfix19_En18 
  input [18:0] Wgt_664, // sfix19_En18 
  input [18:0] Wgt_665, // sfix19_En18 
  input [18:0] Wgt_666, // sfix19_En18 
  input [18:0] Wgt_667, // sfix19_En18 
  input [18:0] Wgt_668, // sfix19_En18 
  input [18:0] Wgt_669, // sfix19_En18 
  input [18:0] Wgt_670, // sfix19_En18 
  input [18:0] Wgt_671, // sfix19_En18 
  input [18:0] Wgt_672, // sfix19_En18 
  input [18:0] Wgt_673, // sfix19_En18 
  input [18:0] Wgt_674, // sfix19_En18 
  input [18:0] Wgt_675, // sfix19_En18 
  input [18:0] Wgt_676, // sfix19_En18 
  input [18:0] Wgt_677, // sfix19_En18 
  input [18:0] Wgt_678, // sfix19_En18 
  input [18:0] Wgt_679, // sfix19_En18 
  input [18:0] Wgt_680, // sfix19_En18 
  input [18:0] Wgt_681, // sfix19_En18 
  input [18:0] Wgt_682, // sfix19_En18 
  input [18:0] Wgt_683, // sfix19_En18 
  input [18:0] Wgt_684, // sfix19_En18 
  input [18:0] Wgt_685, // sfix19_En18 
  input [18:0] Wgt_686, // sfix19_En18 
  input [18:0] Wgt_687, // sfix19_En18 
  input [18:0] Wgt_688, // sfix19_En18 
  input [18:0] Wgt_689, // sfix19_En18 
  input [18:0] Wgt_690, // sfix19_En18 
  input [18:0] Wgt_691, // sfix19_En18 
  input [18:0] Wgt_692, // sfix19_En18 
  input [18:0] Wgt_693, // sfix19_En18 
  input [18:0] Wgt_694, // sfix19_En18 
  input [18:0] Wgt_695, // sfix19_En18 
  input [18:0] Wgt_696, // sfix19_En18 
  input [18:0] Wgt_697, // sfix19_En18 
  input [18:0] Wgt_698, // sfix19_En18 
  input [18:0] Wgt_699, // sfix19_En18 
  input [18:0] Wgt_700, // sfix19_En18 
  input [18:0] Wgt_701, // sfix19_En18 
  input [18:0] Wgt_702, // sfix19_En18 
  input [18:0] Wgt_703, // sfix19_En18 
  input [18:0] Wgt_704, // sfix19_En18 
  input [18:0] Wgt_705, // sfix19_En18 
  input [18:0] Wgt_706, // sfix19_En18 
  input [18:0] Wgt_707, // sfix19_En18 
  input [18:0] Wgt_708, // sfix19_En18 
  input [18:0] Wgt_709, // sfix19_En18 
  input [18:0] Wgt_710, // sfix19_En18 
  input [18:0] Wgt_711, // sfix19_En18 
  input [18:0] Wgt_712, // sfix19_En18 
  input [18:0] Wgt_713, // sfix19_En18 
  input [18:0] Wgt_714, // sfix19_En18 
  input [18:0] Wgt_715, // sfix19_En18 
  input [18:0] Wgt_716, // sfix19_En18 
  input [18:0] Wgt_717, // sfix19_En18 
  input [18:0] Wgt_718, // sfix19_En18 
  input [18:0] Wgt_719, // sfix19_En18 
  input [18:0] Wgt_720, // sfix19_En18 
  input [18:0] Wgt_721, // sfix19_En18 
  input [18:0] Wgt_722, // sfix19_En18 
  input [18:0] Wgt_723, // sfix19_En18 
  input [18:0] Wgt_724, // sfix19_En18 
  input [18:0] Wgt_725, // sfix19_En18 
  input [18:0] Wgt_726, // sfix19_En18 
  input [18:0] Wgt_727, // sfix19_En18 
  input [18:0] Wgt_728, // sfix19_En18 
  input [18:0] Wgt_729, // sfix19_En18 
  input [18:0] Wgt_730, // sfix19_En18 
  input [18:0] Wgt_731, // sfix19_En18 
  input [18:0] Wgt_732, // sfix19_En18 
  input [18:0] Wgt_733, // sfix19_En18 
  input [18:0] Wgt_734, // sfix19_En18 
  input [18:0] Wgt_735, // sfix19_En18 
  input [18:0] Wgt_736, // sfix19_En18 
  input [18:0] Wgt_737, // sfix19_En18 
  input [18:0] Wgt_738, // sfix19_En18 
  input [18:0] Wgt_739, // sfix19_En18 
  input [18:0] Wgt_740, // sfix19_En18 
  input [18:0] Wgt_741, // sfix19_En18 
  input [18:0] Wgt_742, // sfix19_En18 
  input [18:0] Wgt_743, // sfix19_En18 
  input [18:0] Wgt_744, // sfix19_En18 
  input [18:0] Wgt_745, // sfix19_En18 
  input [18:0] Wgt_746, // sfix19_En18 
  input [18:0] Wgt_747, // sfix19_En18 
  input [18:0] Wgt_748, // sfix19_En18 
  input [18:0] Wgt_749, // sfix19_En18 
  input [18:0] Wgt_750, // sfix19_En18 
  input [18:0] Wgt_751, // sfix19_En18 
  input [18:0] Wgt_752, // sfix19_En18 
  input [18:0] Wgt_753, // sfix19_En18 
  input [18:0] Wgt_754, // sfix19_En18 
  input [18:0] Wgt_755, // sfix19_En18 
  input [18:0] Wgt_756, // sfix19_En18 
  input [18:0] Wgt_757, // sfix19_En18 
  input [18:0] Wgt_758, // sfix19_En18 
  input [18:0] Wgt_759, // sfix19_En18 
  input [18:0] Wgt_760, // sfix19_En18 
  input [18:0] Wgt_761, // sfix19_En18 
  input [18:0] Wgt_762, // sfix19_En18 
  input [18:0] Wgt_763, // sfix19_En18 
  input [18:0] Wgt_764, // sfix19_En18 
  input [18:0] Wgt_765, // sfix19_En18 
  input [18:0] Wgt_766, // sfix19_En18 
  input [18:0] Wgt_767, // sfix19_En18 
  input [18:0] Wgt_768, // sfix19_En18 
  input [18:0] Wgt_769, // sfix19_En18 
  input [18:0] Wgt_770, // sfix19_En18 
  input [18:0] Wgt_771, // sfix19_En18 
  input [18:0] Wgt_772, // sfix19_En18 
  input [18:0] Wgt_773, // sfix19_En18 
  input [18:0] Wgt_774, // sfix19_En18 
  input [18:0] Wgt_775, // sfix19_En18 
  input [18:0] Wgt_776, // sfix19_En18 
  input [18:0] Wgt_777, // sfix19_En18 
  input [18:0] Wgt_778, // sfix19_En18 
  input [18:0] Wgt_779, // sfix19_En18 
  input [18:0] Wgt_780, // sfix19_En18 
  input [18:0] Wgt_781, // sfix19_En18 
  input [18:0] Wgt_782, // sfix19_En18 
  input [18:0] Wgt_783, // sfix19_En18 
  input [18:0] Wgt_784, // sfix19_En18 
 output [25:0] cell_out,
 output Output_Valid
	);

reg[5:0] select;
reg [6:0] state;
reg Output_Valid_r;
reg [8:0] counter;
reg [25:0] cell_out_r;
wire [25:0] tot_out;
wire [25:0] tot_out_real;
// 28 outputs, in total the final output
reg [25:0] sum_reg0;
reg [25:0] sum_reg1;
reg [25:0] sum_reg2;
reg [25:0] sum_reg3;
reg [25:0] sum_reg4;
reg [25:0] sum_reg5;
reg [25:0] sum_reg6;
reg [25:0] sum_reg7;
reg [25:0] sum_reg8;
reg [25:0] sum_reg9;
reg [25:0] sum_reg10;
reg [25:0] sum_reg11;
reg [25:0] sum_reg12;
reg [25:0] sum_reg13;
reg [25:0] sum_reg14;
reg [25:0] sum_reg15;
reg [25:0] sum_reg16;
reg [25:0] sum_reg17;
reg [25:0] sum_reg18;
reg [25:0] sum_reg19;
reg [25:0] sum_reg20;
reg [25:0] sum_reg21;
reg [25:0] sum_reg22;
reg [25:0] sum_reg23;
reg [25:0] sum_reg24;
reg [25:0] sum_reg25;
reg [25:0] sum_reg26;
reg [25:0] sum_reg27;


//等28个sum全部出来之后统一赋值统一进入加法器
reg [25:0] sum_sim_reg0;
reg [25:0] sum_sim_reg1;
reg [25:0] sum_sim_reg2;
reg [25:0] sum_sim_reg3;
reg [25:0] sum_sim_reg4;
reg [25:0] sum_sim_reg5;
reg [25:0] sum_sim_reg6;
reg [25:0] sum_sim_reg7;
reg [25:0] sum_sim_reg8;
reg [25:0] sum_sim_reg9;
reg [25:0] sum_sim_reg10;
reg [25:0] sum_sim_reg11;
reg [25:0] sum_sim_reg12;
reg [25:0] sum_sim_reg13;
reg [25:0] sum_sim_reg14;
reg [25:0] sum_sim_reg15;
reg [25:0] sum_sim_reg16;
reg [25:0] sum_sim_reg17;
reg [25:0] sum_sim_reg18;
reg [25:0] sum_sim_reg19;
reg [25:0] sum_sim_reg20;
reg [25:0] sum_sim_reg21;
reg [25:0] sum_sim_reg22;
reg [25:0] sum_sim_reg23;
reg [25:0] sum_sim_reg24;
reg [25:0] sum_sim_reg25;
reg [25:0] sum_sim_reg26;
reg [25:0] sum_sim_reg27;

//所有input全部存一次

reg [9:0] Pix_reg_0;
reg [9:0] Pix_reg_1;
reg [9:0] Pix_reg_2;
reg [9:0] Pix_reg_3;
reg [9:0] Pix_reg_4;
reg [9:0] Pix_reg_5;
reg [9:0] Pix_reg_6;
reg [9:0] Pix_reg_7;
reg [9:0] Pix_reg_8;
reg [9:0] Pix_reg_9;
reg [9:0] Pix_reg_10;
reg [9:0] Pix_reg_11;
reg [9:0] Pix_reg_12;
reg [9:0] Pix_reg_13;
reg [9:0] Pix_reg_14;
reg [9:0] Pix_reg_15;
reg [9:0] Pix_reg_16;
reg [9:0] Pix_reg_17;
reg [9:0] Pix_reg_18;
reg [9:0] Pix_reg_19;
reg [9:0] Pix_reg_20;
reg [9:0] Pix_reg_21;
reg [9:0] Pix_reg_22;
reg [9:0] Pix_reg_23;
reg [9:0] Pix_reg_24;
reg [9:0] Pix_reg_25;
reg [9:0] Pix_reg_26;
reg [9:0] Pix_reg_27;
reg [9:0] Pix_reg_28;
reg [9:0] Pix_reg_29;
reg [9:0] Pix_reg_30;
reg [9:0] Pix_reg_31;
reg [9:0] Pix_reg_32;
reg [9:0] Pix_reg_33;
reg [9:0] Pix_reg_34;
reg [9:0] Pix_reg_35;
reg [9:0] Pix_reg_36;
reg [9:0] Pix_reg_37;
reg [9:0] Pix_reg_38;
reg [9:0] Pix_reg_39;
reg [9:0] Pix_reg_40;
reg [9:0] Pix_reg_41;
reg [9:0] Pix_reg_42;
reg [9:0] Pix_reg_43;
reg [9:0] Pix_reg_44;
reg [9:0] Pix_reg_45;
reg [9:0] Pix_reg_46;
reg [9:0] Pix_reg_47;
reg [9:0] Pix_reg_48;
reg [9:0] Pix_reg_49;
reg [9:0] Pix_reg_50;
reg [9:0] Pix_reg_51;
reg [9:0] Pix_reg_52;
reg [9:0] Pix_reg_53;
reg [9:0] Pix_reg_54;
reg [9:0] Pix_reg_55;
reg [9:0] Pix_reg_56;
reg [9:0] Pix_reg_57;
reg [9:0] Pix_reg_58;
reg [9:0] Pix_reg_59;
reg [9:0] Pix_reg_60;
reg [9:0] Pix_reg_61;
reg [9:0] Pix_reg_62;
reg [9:0] Pix_reg_63;
reg [9:0] Pix_reg_64;
reg [9:0] Pix_reg_65;
reg [9:0] Pix_reg_66;
reg [9:0] Pix_reg_67;
reg [9:0] Pix_reg_68;
reg [9:0] Pix_reg_69;
reg [9:0] Pix_reg_70;
reg [9:0] Pix_reg_71;
reg [9:0] Pix_reg_72;
reg [9:0] Pix_reg_73;
reg [9:0] Pix_reg_74;
reg [9:0] Pix_reg_75;
reg [9:0] Pix_reg_76;
reg [9:0] Pix_reg_77;
reg [9:0] Pix_reg_78;
reg [9:0] Pix_reg_79;
reg [9:0] Pix_reg_80;
reg [9:0] Pix_reg_81;
reg [9:0] Pix_reg_82;
reg [9:0] Pix_reg_83;
reg [9:0] Pix_reg_84;
reg [9:0] Pix_reg_85;
reg [9:0] Pix_reg_86;
reg [9:0] Pix_reg_87;
reg [9:0] Pix_reg_88;
reg [9:0] Pix_reg_89;
reg [9:0] Pix_reg_90;
reg [9:0] Pix_reg_91;
reg [9:0] Pix_reg_92;
reg [9:0] Pix_reg_93;
reg [9:0] Pix_reg_94;
reg [9:0] Pix_reg_95;
reg [9:0] Pix_reg_96;
reg [9:0] Pix_reg_97;
reg [9:0] Pix_reg_98;
reg [9:0] Pix_reg_99;
reg [9:0] Pix_reg_100;
reg [9:0] Pix_reg_101;
reg [9:0] Pix_reg_102;
reg [9:0] Pix_reg_103;
reg [9:0] Pix_reg_104;
reg [9:0] Pix_reg_105;
reg [9:0] Pix_reg_106;
reg [9:0] Pix_reg_107;
reg [9:0] Pix_reg_108;
reg [9:0] Pix_reg_109;
reg [9:0] Pix_reg_110;
reg [9:0] Pix_reg_111;
reg [9:0] Pix_reg_112;
reg [9:0] Pix_reg_113;
reg [9:0] Pix_reg_114;
reg [9:0] Pix_reg_115;
reg [9:0] Pix_reg_116;
reg [9:0] Pix_reg_117;
reg [9:0] Pix_reg_118;
reg [9:0] Pix_reg_119;
reg [9:0] Pix_reg_120;
reg [9:0] Pix_reg_121;
reg [9:0] Pix_reg_122;
reg [9:0] Pix_reg_123;
reg [9:0] Pix_reg_124;
reg [9:0] Pix_reg_125;
reg [9:0] Pix_reg_126;
reg [9:0] Pix_reg_127;
reg [9:0] Pix_reg_128;
reg [9:0] Pix_reg_129;
reg [9:0] Pix_reg_130;
reg [9:0] Pix_reg_131;
reg [9:0] Pix_reg_132;
reg [9:0] Pix_reg_133;
reg [9:0] Pix_reg_134;
reg [9:0] Pix_reg_135;
reg [9:0] Pix_reg_136;
reg [9:0] Pix_reg_137;
reg [9:0] Pix_reg_138;
reg [9:0] Pix_reg_139;
reg [9:0] Pix_reg_140;
reg [9:0] Pix_reg_141;
reg [9:0] Pix_reg_142;
reg [9:0] Pix_reg_143;
reg [9:0] Pix_reg_144;
reg [9:0] Pix_reg_145;
reg [9:0] Pix_reg_146;
reg [9:0] Pix_reg_147;
reg [9:0] Pix_reg_148;
reg [9:0] Pix_reg_149;
reg [9:0] Pix_reg_150;
reg [9:0] Pix_reg_151;
reg [9:0] Pix_reg_152;
reg [9:0] Pix_reg_153;
reg [9:0] Pix_reg_154;
reg [9:0] Pix_reg_155;
reg [9:0] Pix_reg_156;
reg [9:0] Pix_reg_157;
reg [9:0] Pix_reg_158;
reg [9:0] Pix_reg_159;
reg [9:0] Pix_reg_160;
reg [9:0] Pix_reg_161;
reg [9:0] Pix_reg_162;
reg [9:0] Pix_reg_163;
reg [9:0] Pix_reg_164;
reg [9:0] Pix_reg_165;
reg [9:0] Pix_reg_166;
reg [9:0] Pix_reg_167;
reg [9:0] Pix_reg_168;
reg [9:0] Pix_reg_169;
reg [9:0] Pix_reg_170;
reg [9:0] Pix_reg_171;
reg [9:0] Pix_reg_172;
reg [9:0] Pix_reg_173;
reg [9:0] Pix_reg_174;
reg [9:0] Pix_reg_175;
reg [9:0] Pix_reg_176;
reg [9:0] Pix_reg_177;
reg [9:0] Pix_reg_178;
reg [9:0] Pix_reg_179;
reg [9:0] Pix_reg_180;
reg [9:0] Pix_reg_181;
reg [9:0] Pix_reg_182;
reg [9:0] Pix_reg_183;
reg [9:0] Pix_reg_184;
reg [9:0] Pix_reg_185;
reg [9:0] Pix_reg_186;
reg [9:0] Pix_reg_187;
reg [9:0] Pix_reg_188;
reg [9:0] Pix_reg_189;
reg [9:0] Pix_reg_190;
reg [9:0] Pix_reg_191;
reg [9:0] Pix_reg_192;
reg [9:0] Pix_reg_193;
reg [9:0] Pix_reg_194;
reg [9:0] Pix_reg_195;
reg [9:0] Pix_reg_196;
reg [9:0] Pix_reg_197;
reg [9:0] Pix_reg_198;
reg [9:0] Pix_reg_199;
reg [9:0] Pix_reg_200;
reg [9:0] Pix_reg_201;
reg [9:0] Pix_reg_202;
reg [9:0] Pix_reg_203;
reg [9:0] Pix_reg_204;
reg [9:0] Pix_reg_205;
reg [9:0] Pix_reg_206;
reg [9:0] Pix_reg_207;
reg [9:0] Pix_reg_208;
reg [9:0] Pix_reg_209;
reg [9:0] Pix_reg_210;
reg [9:0] Pix_reg_211;
reg [9:0] Pix_reg_212;
reg [9:0] Pix_reg_213;
reg [9:0] Pix_reg_214;
reg [9:0] Pix_reg_215;
reg [9:0] Pix_reg_216;
reg [9:0] Pix_reg_217;
reg [9:0] Pix_reg_218;
reg [9:0] Pix_reg_219;
reg [9:0] Pix_reg_220;
reg [9:0] Pix_reg_221;
reg [9:0] Pix_reg_222;
reg [9:0] Pix_reg_223;
reg [9:0] Pix_reg_224;
reg [9:0] Pix_reg_225;
reg [9:0] Pix_reg_226;
reg [9:0] Pix_reg_227;
reg [9:0] Pix_reg_228;
reg [9:0] Pix_reg_229;
reg [9:0] Pix_reg_230;
reg [9:0] Pix_reg_231;
reg [9:0] Pix_reg_232;
reg [9:0] Pix_reg_233;
reg [9:0] Pix_reg_234;
reg [9:0] Pix_reg_235;
reg [9:0] Pix_reg_236;
reg [9:0] Pix_reg_237;
reg [9:0] Pix_reg_238;
reg [9:0] Pix_reg_239;
reg [9:0] Pix_reg_240;
reg [9:0] Pix_reg_241;
reg [9:0] Pix_reg_242;
reg [9:0] Pix_reg_243;
reg [9:0] Pix_reg_244;
reg [9:0] Pix_reg_245;
reg [9:0] Pix_reg_246;
reg [9:0] Pix_reg_247;
reg [9:0] Pix_reg_248;
reg [9:0] Pix_reg_249;
reg [9:0] Pix_reg_250;
reg [9:0] Pix_reg_251;
reg [9:0] Pix_reg_252;
reg [9:0] Pix_reg_253;
reg [9:0] Pix_reg_254;
reg [9:0] Pix_reg_255;
reg [9:0] Pix_reg_256;
reg [9:0] Pix_reg_257;
reg [9:0] Pix_reg_258;
reg [9:0] Pix_reg_259;
reg [9:0] Pix_reg_260;
reg [9:0] Pix_reg_261;
reg [9:0] Pix_reg_262;
reg [9:0] Pix_reg_263;
reg [9:0] Pix_reg_264;
reg [9:0] Pix_reg_265;
reg [9:0] Pix_reg_266;
reg [9:0] Pix_reg_267;
reg [9:0] Pix_reg_268;
reg [9:0] Pix_reg_269;
reg [9:0] Pix_reg_270;
reg [9:0] Pix_reg_271;
reg [9:0] Pix_reg_272;
reg [9:0] Pix_reg_273;
reg [9:0] Pix_reg_274;
reg [9:0] Pix_reg_275;
reg [9:0] Pix_reg_276;
reg [9:0] Pix_reg_277;
reg [9:0] Pix_reg_278;
reg [9:0] Pix_reg_279;
reg [9:0] Pix_reg_280;
reg [9:0] Pix_reg_281;
reg [9:0] Pix_reg_282;
reg [9:0] Pix_reg_283;
reg [9:0] Pix_reg_284;
reg [9:0] Pix_reg_285;
reg [9:0] Pix_reg_286;
reg [9:0] Pix_reg_287;
reg [9:0] Pix_reg_288;
reg [9:0] Pix_reg_289;
reg [9:0] Pix_reg_290;
reg [9:0] Pix_reg_291;
reg [9:0] Pix_reg_292;
reg [9:0] Pix_reg_293;
reg [9:0] Pix_reg_294;
reg [9:0] Pix_reg_295;
reg [9:0] Pix_reg_296;
reg [9:0] Pix_reg_297;
reg [9:0] Pix_reg_298;
reg [9:0] Pix_reg_299;
reg [9:0] Pix_reg_300;
reg [9:0] Pix_reg_301;
reg [9:0] Pix_reg_302;
reg [9:0] Pix_reg_303;
reg [9:0] Pix_reg_304;
reg [9:0] Pix_reg_305;
reg [9:0] Pix_reg_306;
reg [9:0] Pix_reg_307;
reg [9:0] Pix_reg_308;
reg [9:0] Pix_reg_309;
reg [9:0] Pix_reg_310;
reg [9:0] Pix_reg_311;
reg [9:0] Pix_reg_312;
reg [9:0] Pix_reg_313;
reg [9:0] Pix_reg_314;
reg [9:0] Pix_reg_315;
reg [9:0] Pix_reg_316;
reg [9:0] Pix_reg_317;
reg [9:0] Pix_reg_318;
reg [9:0] Pix_reg_319;
reg [9:0] Pix_reg_320;
reg [9:0] Pix_reg_321;
reg [9:0] Pix_reg_322;
reg [9:0] Pix_reg_323;
reg [9:0] Pix_reg_324;
reg [9:0] Pix_reg_325;
reg [9:0] Pix_reg_326;
reg [9:0] Pix_reg_327;
reg [9:0] Pix_reg_328;
reg [9:0] Pix_reg_329;
reg [9:0] Pix_reg_330;
reg [9:0] Pix_reg_331;
reg [9:0] Pix_reg_332;
reg [9:0] Pix_reg_333;
reg [9:0] Pix_reg_334;
reg [9:0] Pix_reg_335;
reg [9:0] Pix_reg_336;
reg [9:0] Pix_reg_337;
reg [9:0] Pix_reg_338;
reg [9:0] Pix_reg_339;
reg [9:0] Pix_reg_340;
reg [9:0] Pix_reg_341;
reg [9:0] Pix_reg_342;
reg [9:0] Pix_reg_343;
reg [9:0] Pix_reg_344;
reg [9:0] Pix_reg_345;
reg [9:0] Pix_reg_346;
reg [9:0] Pix_reg_347;
reg [9:0] Pix_reg_348;
reg [9:0] Pix_reg_349;
reg [9:0] Pix_reg_350;
reg [9:0] Pix_reg_351;
reg [9:0] Pix_reg_352;
reg [9:0] Pix_reg_353;
reg [9:0] Pix_reg_354;
reg [9:0] Pix_reg_355;
reg [9:0] Pix_reg_356;
reg [9:0] Pix_reg_357;
reg [9:0] Pix_reg_358;
reg [9:0] Pix_reg_359;
reg [9:0] Pix_reg_360;
reg [9:0] Pix_reg_361;
reg [9:0] Pix_reg_362;
reg [9:0] Pix_reg_363;
reg [9:0] Pix_reg_364;
reg [9:0] Pix_reg_365;
reg [9:0] Pix_reg_366;
reg [9:0] Pix_reg_367;
reg [9:0] Pix_reg_368;
reg [9:0] Pix_reg_369;
reg [9:0] Pix_reg_370;
reg [9:0] Pix_reg_371;
reg [9:0] Pix_reg_372;
reg [9:0] Pix_reg_373;
reg [9:0] Pix_reg_374;
reg [9:0] Pix_reg_375;
reg [9:0] Pix_reg_376;
reg [9:0] Pix_reg_377;
reg [9:0] Pix_reg_378;
reg [9:0] Pix_reg_379;
reg [9:0] Pix_reg_380;
reg [9:0] Pix_reg_381;
reg [9:0] Pix_reg_382;
reg [9:0] Pix_reg_383;
reg [9:0] Pix_reg_384;
reg [9:0] Pix_reg_385;
reg [9:0] Pix_reg_386;
reg [9:0] Pix_reg_387;
reg [9:0] Pix_reg_388;
reg [9:0] Pix_reg_389;
reg [9:0] Pix_reg_390;
reg [9:0] Pix_reg_391;
reg [9:0] Pix_reg_392;
reg [9:0] Pix_reg_393;
reg [9:0] Pix_reg_394;
reg [9:0] Pix_reg_395;
reg [9:0] Pix_reg_396;
reg [9:0] Pix_reg_397;
reg [9:0] Pix_reg_398;
reg [9:0] Pix_reg_399;
reg [9:0] Pix_reg_400;
reg [9:0] Pix_reg_401;
reg [9:0] Pix_reg_402;
reg [9:0] Pix_reg_403;
reg [9:0] Pix_reg_404;
reg [9:0] Pix_reg_405;
reg [9:0] Pix_reg_406;
reg [9:0] Pix_reg_407;
reg [9:0] Pix_reg_408;
reg [9:0] Pix_reg_409;
reg [9:0] Pix_reg_410;
reg [9:0] Pix_reg_411;
reg [9:0] Pix_reg_412;
reg [9:0] Pix_reg_413;
reg [9:0] Pix_reg_414;
reg [9:0] Pix_reg_415;
reg [9:0] Pix_reg_416;
reg [9:0] Pix_reg_417;
reg [9:0] Pix_reg_418;
reg [9:0] Pix_reg_419;
reg [9:0] Pix_reg_420;
reg [9:0] Pix_reg_421;
reg [9:0] Pix_reg_422;
reg [9:0] Pix_reg_423;
reg [9:0] Pix_reg_424;
reg [9:0] Pix_reg_425;
reg [9:0] Pix_reg_426;
reg [9:0] Pix_reg_427;
reg [9:0] Pix_reg_428;
reg [9:0] Pix_reg_429;
reg [9:0] Pix_reg_430;
reg [9:0] Pix_reg_431;
reg [9:0] Pix_reg_432;
reg [9:0] Pix_reg_433;
reg [9:0] Pix_reg_434;
reg [9:0] Pix_reg_435;
reg [9:0] Pix_reg_436;
reg [9:0] Pix_reg_437;
reg [9:0] Pix_reg_438;
reg [9:0] Pix_reg_439;
reg [9:0] Pix_reg_440;
reg [9:0] Pix_reg_441;
reg [9:0] Pix_reg_442;
reg [9:0] Pix_reg_443;
reg [9:0] Pix_reg_444;
reg [9:0] Pix_reg_445;
reg [9:0] Pix_reg_446;
reg [9:0] Pix_reg_447;
reg [9:0] Pix_reg_448;
reg [9:0] Pix_reg_449;
reg [9:0] Pix_reg_450;
reg [9:0] Pix_reg_451;
reg [9:0] Pix_reg_452;
reg [9:0] Pix_reg_453;
reg [9:0] Pix_reg_454;
reg [9:0] Pix_reg_455;
reg [9:0] Pix_reg_456;
reg [9:0] Pix_reg_457;
reg [9:0] Pix_reg_458;
reg [9:0] Pix_reg_459;
reg [9:0] Pix_reg_460;
reg [9:0] Pix_reg_461;
reg [9:0] Pix_reg_462;
reg [9:0] Pix_reg_463;
reg [9:0] Pix_reg_464;
reg [9:0] Pix_reg_465;
reg [9:0] Pix_reg_466;
reg [9:0] Pix_reg_467;
reg [9:0] Pix_reg_468;
reg [9:0] Pix_reg_469;
reg [9:0] Pix_reg_470;
reg [9:0] Pix_reg_471;
reg [9:0] Pix_reg_472;
reg [9:0] Pix_reg_473;
reg [9:0] Pix_reg_474;
reg [9:0] Pix_reg_475;
reg [9:0] Pix_reg_476;
reg [9:0] Pix_reg_477;
reg [9:0] Pix_reg_478;
reg [9:0] Pix_reg_479;
reg [9:0] Pix_reg_480;
reg [9:0] Pix_reg_481;
reg [9:0] Pix_reg_482;
reg [9:0] Pix_reg_483;
reg [9:0] Pix_reg_484;
reg [9:0] Pix_reg_485;
reg [9:0] Pix_reg_486;
reg [9:0] Pix_reg_487;
reg [9:0] Pix_reg_488;
reg [9:0] Pix_reg_489;
reg [9:0] Pix_reg_490;
reg [9:0] Pix_reg_491;
reg [9:0] Pix_reg_492;
reg [9:0] Pix_reg_493;
reg [9:0] Pix_reg_494;
reg [9:0] Pix_reg_495;
reg [9:0] Pix_reg_496;
reg [9:0] Pix_reg_497;
reg [9:0] Pix_reg_498;
reg [9:0] Pix_reg_499;
reg [9:0] Pix_reg_500;
reg [9:0] Pix_reg_501;
reg [9:0] Pix_reg_502;
reg [9:0] Pix_reg_503;
reg [9:0] Pix_reg_504;
reg [9:0] Pix_reg_505;
reg [9:0] Pix_reg_506;
reg [9:0] Pix_reg_507;
reg [9:0] Pix_reg_508;
reg [9:0] Pix_reg_509;
reg [9:0] Pix_reg_510;
reg [9:0] Pix_reg_511;
reg [9:0] Pix_reg_512;
reg [9:0] Pix_reg_513;
reg [9:0] Pix_reg_514;
reg [9:0] Pix_reg_515;
reg [9:0] Pix_reg_516;
reg [9:0] Pix_reg_517;
reg [9:0] Pix_reg_518;
reg [9:0] Pix_reg_519;
reg [9:0] Pix_reg_520;
reg [9:0] Pix_reg_521;
reg [9:0] Pix_reg_522;
reg [9:0] Pix_reg_523;
reg [9:0] Pix_reg_524;
reg [9:0] Pix_reg_525;
reg [9:0] Pix_reg_526;
reg [9:0] Pix_reg_527;
reg [9:0] Pix_reg_528;
reg [9:0] Pix_reg_529;
reg [9:0] Pix_reg_530;
reg [9:0] Pix_reg_531;
reg [9:0] Pix_reg_532;
reg [9:0] Pix_reg_533;
reg [9:0] Pix_reg_534;
reg [9:0] Pix_reg_535;
reg [9:0] Pix_reg_536;
reg [9:0] Pix_reg_537;
reg [9:0] Pix_reg_538;
reg [9:0] Pix_reg_539;
reg [9:0] Pix_reg_540;
reg [9:0] Pix_reg_541;
reg [9:0] Pix_reg_542;
reg [9:0] Pix_reg_543;
reg [9:0] Pix_reg_544;
reg [9:0] Pix_reg_545;
reg [9:0] Pix_reg_546;
reg [9:0] Pix_reg_547;
reg [9:0] Pix_reg_548;
reg [9:0] Pix_reg_549;
reg [9:0] Pix_reg_550;
reg [9:0] Pix_reg_551;
reg [9:0] Pix_reg_552;
reg [9:0] Pix_reg_553;
reg [9:0] Pix_reg_554;
reg [9:0] Pix_reg_555;
reg [9:0] Pix_reg_556;
reg [9:0] Pix_reg_557;
reg [9:0] Pix_reg_558;
reg [9:0] Pix_reg_559;
reg [9:0] Pix_reg_560;
reg [9:0] Pix_reg_561;
reg [9:0] Pix_reg_562;
reg [9:0] Pix_reg_563;
reg [9:0] Pix_reg_564;
reg [9:0] Pix_reg_565;
reg [9:0] Pix_reg_566;
reg [9:0] Pix_reg_567;
reg [9:0] Pix_reg_568;
reg [9:0] Pix_reg_569;
reg [9:0] Pix_reg_570;
reg [9:0] Pix_reg_571;
reg [9:0] Pix_reg_572;
reg [9:0] Pix_reg_573;
reg [9:0] Pix_reg_574;
reg [9:0] Pix_reg_575;
reg [9:0] Pix_reg_576;
reg [9:0] Pix_reg_577;
reg [9:0] Pix_reg_578;
reg [9:0] Pix_reg_579;
reg [9:0] Pix_reg_580;
reg [9:0] Pix_reg_581;
reg [9:0] Pix_reg_582;
reg [9:0] Pix_reg_583;
reg [9:0] Pix_reg_584;
reg [9:0] Pix_reg_585;
reg [9:0] Pix_reg_586;
reg [9:0] Pix_reg_587;
reg [9:0] Pix_reg_588;
reg [9:0] Pix_reg_589;
reg [9:0] Pix_reg_590;
reg [9:0] Pix_reg_591;
reg [9:0] Pix_reg_592;
reg [9:0] Pix_reg_593;
reg [9:0] Pix_reg_594;
reg [9:0] Pix_reg_595;
reg [9:0] Pix_reg_596;
reg [9:0] Pix_reg_597;
reg [9:0] Pix_reg_598;
reg [9:0] Pix_reg_599;
reg [9:0] Pix_reg_600;
reg [9:0] Pix_reg_601;
reg [9:0] Pix_reg_602;
reg [9:0] Pix_reg_603;
reg [9:0] Pix_reg_604;
reg [9:0] Pix_reg_605;
reg [9:0] Pix_reg_606;
reg [9:0] Pix_reg_607;
reg [9:0] Pix_reg_608;
reg [9:0] Pix_reg_609;
reg [9:0] Pix_reg_610;
reg [9:0] Pix_reg_611;
reg [9:0] Pix_reg_612;
reg [9:0] Pix_reg_613;
reg [9:0] Pix_reg_614;
reg [9:0] Pix_reg_615;
reg [9:0] Pix_reg_616;
reg [9:0] Pix_reg_617;
reg [9:0] Pix_reg_618;
reg [9:0] Pix_reg_619;
reg [9:0] Pix_reg_620;
reg [9:0] Pix_reg_621;
reg [9:0] Pix_reg_622;
reg [9:0] Pix_reg_623;
reg [9:0] Pix_reg_624;
reg [9:0] Pix_reg_625;
reg [9:0] Pix_reg_626;
reg [9:0] Pix_reg_627;
reg [9:0] Pix_reg_628;
reg [9:0] Pix_reg_629;
reg [9:0] Pix_reg_630;
reg [9:0] Pix_reg_631;
reg [9:0] Pix_reg_632;
reg [9:0] Pix_reg_633;
reg [9:0] Pix_reg_634;
reg [9:0] Pix_reg_635;
reg [9:0] Pix_reg_636;
reg [9:0] Pix_reg_637;
reg [9:0] Pix_reg_638;
reg [9:0] Pix_reg_639;
reg [9:0] Pix_reg_640;
reg [9:0] Pix_reg_641;
reg [9:0] Pix_reg_642;
reg [9:0] Pix_reg_643;
reg [9:0] Pix_reg_644;
reg [9:0] Pix_reg_645;
reg [9:0] Pix_reg_646;
reg [9:0] Pix_reg_647;
reg [9:0] Pix_reg_648;
reg [9:0] Pix_reg_649;
reg [9:0] Pix_reg_650;
reg [9:0] Pix_reg_651;
reg [9:0] Pix_reg_652;
reg [9:0] Pix_reg_653;
reg [9:0] Pix_reg_654;
reg [9:0] Pix_reg_655;
reg [9:0] Pix_reg_656;
reg [9:0] Pix_reg_657;
reg [9:0] Pix_reg_658;
reg [9:0] Pix_reg_659;
reg [9:0] Pix_reg_660;
reg [9:0] Pix_reg_661;
reg [9:0] Pix_reg_662;
reg [9:0] Pix_reg_663;
reg [9:0] Pix_reg_664;
reg [9:0] Pix_reg_665;
reg [9:0] Pix_reg_666;
reg [9:0] Pix_reg_667;
reg [9:0] Pix_reg_668;
reg [9:0] Pix_reg_669;
reg [9:0] Pix_reg_670;
reg [9:0] Pix_reg_671;
reg [9:0] Pix_reg_672;
reg [9:0] Pix_reg_673;
reg [9:0] Pix_reg_674;
reg [9:0] Pix_reg_675;
reg [9:0] Pix_reg_676;
reg [9:0] Pix_reg_677;
reg [9:0] Pix_reg_678;
reg [9:0] Pix_reg_679;
reg [9:0] Pix_reg_680;
reg [9:0] Pix_reg_681;
reg [9:0] Pix_reg_682;
reg [9:0] Pix_reg_683;
reg [9:0] Pix_reg_684;
reg [9:0] Pix_reg_685;
reg [9:0] Pix_reg_686;
reg [9:0] Pix_reg_687;
reg [9:0] Pix_reg_688;
reg [9:0] Pix_reg_689;
reg [9:0] Pix_reg_690;
reg [9:0] Pix_reg_691;
reg [9:0] Pix_reg_692;
reg [9:0] Pix_reg_693;
reg [9:0] Pix_reg_694;
reg [9:0] Pix_reg_695;
reg [9:0] Pix_reg_696;
reg [9:0] Pix_reg_697;
reg [9:0] Pix_reg_698;
reg [9:0] Pix_reg_699;
reg [9:0] Pix_reg_700;
reg [9:0] Pix_reg_701;
reg [9:0] Pix_reg_702;
reg [9:0] Pix_reg_703;
reg [9:0] Pix_reg_704;
reg [9:0] Pix_reg_705;
reg [9:0] Pix_reg_706;
reg [9:0] Pix_reg_707;
reg [9:0] Pix_reg_708;
reg [9:0] Pix_reg_709;
reg [9:0] Pix_reg_710;
reg [9:0] Pix_reg_711;
reg [9:0] Pix_reg_712;
reg [9:0] Pix_reg_713;
reg [9:0] Pix_reg_714;
reg [9:0] Pix_reg_715;
reg [9:0] Pix_reg_716;
reg [9:0] Pix_reg_717;
reg [9:0] Pix_reg_718;
reg [9:0] Pix_reg_719;
reg [9:0] Pix_reg_720;
reg [9:0] Pix_reg_721;
reg [9:0] Pix_reg_722;
reg [9:0] Pix_reg_723;
reg [9:0] Pix_reg_724;
reg [9:0] Pix_reg_725;
reg [9:0] Pix_reg_726;
reg [9:0] Pix_reg_727;
reg [9:0] Pix_reg_728;
reg [9:0] Pix_reg_729;
reg [9:0] Pix_reg_730;
reg [9:0] Pix_reg_731;
reg [9:0] Pix_reg_732;
reg [9:0] Pix_reg_733;
reg [9:0] Pix_reg_734;
reg [9:0] Pix_reg_735;
reg [9:0] Pix_reg_736;
reg [9:0] Pix_reg_737;
reg [9:0] Pix_reg_738;
reg [9:0] Pix_reg_739;
reg [9:0] Pix_reg_740;
reg [9:0] Pix_reg_741;
reg [9:0] Pix_reg_742;
reg [9:0] Pix_reg_743;
reg [9:0] Pix_reg_744;
reg [9:0] Pix_reg_745;
reg [9:0] Pix_reg_746;
reg [9:0] Pix_reg_747;
reg [9:0] Pix_reg_748;
reg [9:0] Pix_reg_749;
reg [9:0] Pix_reg_750;
reg [9:0] Pix_reg_751;
reg [9:0] Pix_reg_752;
reg [9:0] Pix_reg_753;
reg [9:0] Pix_reg_754;
reg [9:0] Pix_reg_755;
reg [9:0] Pix_reg_756;
reg [9:0] Pix_reg_757;
reg [9:0] Pix_reg_758;
reg [9:0] Pix_reg_759;
reg [9:0] Pix_reg_760;
reg [9:0] Pix_reg_761;
reg [9:0] Pix_reg_762;
reg [9:0] Pix_reg_763;
reg [9:0] Pix_reg_764;
reg [9:0] Pix_reg_765;
reg [9:0] Pix_reg_766;
reg [9:0] Pix_reg_767;
reg [9:0] Pix_reg_768;
reg [9:0] Pix_reg_769;
reg [9:0] Pix_reg_770;
reg [9:0] Pix_reg_771;
reg [9:0] Pix_reg_772;
reg [9:0] Pix_reg_773;
reg [9:0] Pix_reg_774;
reg [9:0] Pix_reg_775;
reg [9:0] Pix_reg_776;
reg [9:0] Pix_reg_777;
reg [9:0] Pix_reg_778;
reg [9:0] Pix_reg_779;
reg [9:0] Pix_reg_780;
reg [9:0] Pix_reg_781;
reg [9:0] Pix_reg_782;
reg [9:0] Pix_reg_783;
reg [9:0] Pix_reg_784;

reg [18:0] Wgt_reg_0;
reg [18:0] Wgt_reg_1;
reg [18:0] Wgt_reg_2;
reg [18:0] Wgt_reg_3;
reg [18:0] Wgt_reg_4;
reg [18:0] Wgt_reg_5;
reg [18:0] Wgt_reg_6;
reg [18:0] Wgt_reg_7;
reg [18:0] Wgt_reg_8;
reg [18:0] Wgt_reg_9;
reg [18:0] Wgt_reg_10;
reg [18:0] Wgt_reg_11;
reg [18:0] Wgt_reg_12;
reg [18:0] Wgt_reg_13;
reg [18:0] Wgt_reg_14;
reg [18:0] Wgt_reg_15;
reg [18:0] Wgt_reg_16;
reg [18:0] Wgt_reg_17;
reg [18:0] Wgt_reg_18;
reg [18:0] Wgt_reg_19;
reg [18:0] Wgt_reg_20;
reg [18:0] Wgt_reg_21;
reg [18:0] Wgt_reg_22;
reg [18:0] Wgt_reg_23;
reg [18:0] Wgt_reg_24;
reg [18:0] Wgt_reg_25;
reg [18:0] Wgt_reg_26;
reg [18:0] Wgt_reg_27;
reg [18:0] Wgt_reg_28;
reg [18:0] Wgt_reg_29;
reg [18:0] Wgt_reg_30;
reg [18:0] Wgt_reg_31;
reg [18:0] Wgt_reg_32;
reg [18:0] Wgt_reg_33;
reg [18:0] Wgt_reg_34;
reg [18:0] Wgt_reg_35;
reg [18:0] Wgt_reg_36;
reg [18:0] Wgt_reg_37;
reg [18:0] Wgt_reg_38;
reg [18:0] Wgt_reg_39;
reg [18:0] Wgt_reg_40;
reg [18:0] Wgt_reg_41;
reg [18:0] Wgt_reg_42;
reg [18:0] Wgt_reg_43;
reg [18:0] Wgt_reg_44;
reg [18:0] Wgt_reg_45;
reg [18:0] Wgt_reg_46;
reg [18:0] Wgt_reg_47;
reg [18:0] Wgt_reg_48;
reg [18:0] Wgt_reg_49;
reg [18:0] Wgt_reg_50;
reg [18:0] Wgt_reg_51;
reg [18:0] Wgt_reg_52;
reg [18:0] Wgt_reg_53;
reg [18:0] Wgt_reg_54;
reg [18:0] Wgt_reg_55;
reg [18:0] Wgt_reg_56;
reg [18:0] Wgt_reg_57;
reg [18:0] Wgt_reg_58;
reg [18:0] Wgt_reg_59;
reg [18:0] Wgt_reg_60;
reg [18:0] Wgt_reg_61;
reg [18:0] Wgt_reg_62;
reg [18:0] Wgt_reg_63;
reg [18:0] Wgt_reg_64;
reg [18:0] Wgt_reg_65;
reg [18:0] Wgt_reg_66;
reg [18:0] Wgt_reg_67;
reg [18:0] Wgt_reg_68;
reg [18:0] Wgt_reg_69;
reg [18:0] Wgt_reg_70;
reg [18:0] Wgt_reg_71;
reg [18:0] Wgt_reg_72;
reg [18:0] Wgt_reg_73;
reg [18:0] Wgt_reg_74;
reg [18:0] Wgt_reg_75;
reg [18:0] Wgt_reg_76;
reg [18:0] Wgt_reg_77;
reg [18:0] Wgt_reg_78;
reg [18:0] Wgt_reg_79;
reg [18:0] Wgt_reg_80;
reg [18:0] Wgt_reg_81;
reg [18:0] Wgt_reg_82;
reg [18:0] Wgt_reg_83;
reg [18:0] Wgt_reg_84;
reg [18:0] Wgt_reg_85;
reg [18:0] Wgt_reg_86;
reg [18:0] Wgt_reg_87;
reg [18:0] Wgt_reg_88;
reg [18:0] Wgt_reg_89;
reg [18:0] Wgt_reg_90;
reg [18:0] Wgt_reg_91;
reg [18:0] Wgt_reg_92;
reg [18:0] Wgt_reg_93;
reg [18:0] Wgt_reg_94;
reg [18:0] Wgt_reg_95;
reg [18:0] Wgt_reg_96;
reg [18:0] Wgt_reg_97;
reg [18:0] Wgt_reg_98;
reg [18:0] Wgt_reg_99;
reg [18:0] Wgt_reg_100;
reg [18:0] Wgt_reg_101;
reg [18:0] Wgt_reg_102;
reg [18:0] Wgt_reg_103;
reg [18:0] Wgt_reg_104;
reg [18:0] Wgt_reg_105;
reg [18:0] Wgt_reg_106;
reg [18:0] Wgt_reg_107;
reg [18:0] Wgt_reg_108;
reg [18:0] Wgt_reg_109;
reg [18:0] Wgt_reg_110;
reg [18:0] Wgt_reg_111;
reg [18:0] Wgt_reg_112;
reg [18:0] Wgt_reg_113;
reg [18:0] Wgt_reg_114;
reg [18:0] Wgt_reg_115;
reg [18:0] Wgt_reg_116;
reg [18:0] Wgt_reg_117;
reg [18:0] Wgt_reg_118;
reg [18:0] Wgt_reg_119;
reg [18:0] Wgt_reg_120;
reg [18:0] Wgt_reg_121;
reg [18:0] Wgt_reg_122;
reg [18:0] Wgt_reg_123;
reg [18:0] Wgt_reg_124;
reg [18:0] Wgt_reg_125;
reg [18:0] Wgt_reg_126;
reg [18:0] Wgt_reg_127;
reg [18:0] Wgt_reg_128;
reg [18:0] Wgt_reg_129;
reg [18:0] Wgt_reg_130;
reg [18:0] Wgt_reg_131;
reg [18:0] Wgt_reg_132;
reg [18:0] Wgt_reg_133;
reg [18:0] Wgt_reg_134;
reg [18:0] Wgt_reg_135;
reg [18:0] Wgt_reg_136;
reg [18:0] Wgt_reg_137;
reg [18:0] Wgt_reg_138;
reg [18:0] Wgt_reg_139;
reg [18:0] Wgt_reg_140;
reg [18:0] Wgt_reg_141;
reg [18:0] Wgt_reg_142;
reg [18:0] Wgt_reg_143;
reg [18:0] Wgt_reg_144;
reg [18:0] Wgt_reg_145;
reg [18:0] Wgt_reg_146;
reg [18:0] Wgt_reg_147;
reg [18:0] Wgt_reg_148;
reg [18:0] Wgt_reg_149;
reg [18:0] Wgt_reg_150;
reg [18:0] Wgt_reg_151;
reg [18:0] Wgt_reg_152;
reg [18:0] Wgt_reg_153;
reg [18:0] Wgt_reg_154;
reg [18:0] Wgt_reg_155;
reg [18:0] Wgt_reg_156;
reg [18:0] Wgt_reg_157;
reg [18:0] Wgt_reg_158;
reg [18:0] Wgt_reg_159;
reg [18:0] Wgt_reg_160;
reg [18:0] Wgt_reg_161;
reg [18:0] Wgt_reg_162;
reg [18:0] Wgt_reg_163;
reg [18:0] Wgt_reg_164;
reg [18:0] Wgt_reg_165;
reg [18:0] Wgt_reg_166;
reg [18:0] Wgt_reg_167;
reg [18:0] Wgt_reg_168;
reg [18:0] Wgt_reg_169;
reg [18:0] Wgt_reg_170;
reg [18:0] Wgt_reg_171;
reg [18:0] Wgt_reg_172;
reg [18:0] Wgt_reg_173;
reg [18:0] Wgt_reg_174;
reg [18:0] Wgt_reg_175;
reg [18:0] Wgt_reg_176;
reg [18:0] Wgt_reg_177;
reg [18:0] Wgt_reg_178;
reg [18:0] Wgt_reg_179;
reg [18:0] Wgt_reg_180;
reg [18:0] Wgt_reg_181;
reg [18:0] Wgt_reg_182;
reg [18:0] Wgt_reg_183;
reg [18:0] Wgt_reg_184;
reg [18:0] Wgt_reg_185;
reg [18:0] Wgt_reg_186;
reg [18:0] Wgt_reg_187;
reg [18:0] Wgt_reg_188;
reg [18:0] Wgt_reg_189;
reg [18:0] Wgt_reg_190;
reg [18:0] Wgt_reg_191;
reg [18:0] Wgt_reg_192;
reg [18:0] Wgt_reg_193;
reg [18:0] Wgt_reg_194;
reg [18:0] Wgt_reg_195;
reg [18:0] Wgt_reg_196;
reg [18:0] Wgt_reg_197;
reg [18:0] Wgt_reg_198;
reg [18:0] Wgt_reg_199;
reg [18:0] Wgt_reg_200;
reg [18:0] Wgt_reg_201;
reg [18:0] Wgt_reg_202;
reg [18:0] Wgt_reg_203;
reg [18:0] Wgt_reg_204;
reg [18:0] Wgt_reg_205;
reg [18:0] Wgt_reg_206;
reg [18:0] Wgt_reg_207;
reg [18:0] Wgt_reg_208;
reg [18:0] Wgt_reg_209;
reg [18:0] Wgt_reg_210;
reg [18:0] Wgt_reg_211;
reg [18:0] Wgt_reg_212;
reg [18:0] Wgt_reg_213;
reg [18:0] Wgt_reg_214;
reg [18:0] Wgt_reg_215;
reg [18:0] Wgt_reg_216;
reg [18:0] Wgt_reg_217;
reg [18:0] Wgt_reg_218;
reg [18:0] Wgt_reg_219;
reg [18:0] Wgt_reg_220;
reg [18:0] Wgt_reg_221;
reg [18:0] Wgt_reg_222;
reg [18:0] Wgt_reg_223;
reg [18:0] Wgt_reg_224;
reg [18:0] Wgt_reg_225;
reg [18:0] Wgt_reg_226;
reg [18:0] Wgt_reg_227;
reg [18:0] Wgt_reg_228;
reg [18:0] Wgt_reg_229;
reg [18:0] Wgt_reg_230;
reg [18:0] Wgt_reg_231;
reg [18:0] Wgt_reg_232;
reg [18:0] Wgt_reg_233;
reg [18:0] Wgt_reg_234;
reg [18:0] Wgt_reg_235;
reg [18:0] Wgt_reg_236;
reg [18:0] Wgt_reg_237;
reg [18:0] Wgt_reg_238;
reg [18:0] Wgt_reg_239;
reg [18:0] Wgt_reg_240;
reg [18:0] Wgt_reg_241;
reg [18:0] Wgt_reg_242;
reg [18:0] Wgt_reg_243;
reg [18:0] Wgt_reg_244;
reg [18:0] Wgt_reg_245;
reg [18:0] Wgt_reg_246;
reg [18:0] Wgt_reg_247;
reg [18:0] Wgt_reg_248;
reg [18:0] Wgt_reg_249;
reg [18:0] Wgt_reg_250;
reg [18:0] Wgt_reg_251;
reg [18:0] Wgt_reg_252;
reg [18:0] Wgt_reg_253;
reg [18:0] Wgt_reg_254;
reg [18:0] Wgt_reg_255;
reg [18:0] Wgt_reg_256;
reg [18:0] Wgt_reg_257;
reg [18:0] Wgt_reg_258;
reg [18:0] Wgt_reg_259;
reg [18:0] Wgt_reg_260;
reg [18:0] Wgt_reg_261;
reg [18:0] Wgt_reg_262;
reg [18:0] Wgt_reg_263;
reg [18:0] Wgt_reg_264;
reg [18:0] Wgt_reg_265;
reg [18:0] Wgt_reg_266;
reg [18:0] Wgt_reg_267;
reg [18:0] Wgt_reg_268;
reg [18:0] Wgt_reg_269;
reg [18:0] Wgt_reg_270;
reg [18:0] Wgt_reg_271;
reg [18:0] Wgt_reg_272;
reg [18:0] Wgt_reg_273;
reg [18:0] Wgt_reg_274;
reg [18:0] Wgt_reg_275;
reg [18:0] Wgt_reg_276;
reg [18:0] Wgt_reg_277;
reg [18:0] Wgt_reg_278;
reg [18:0] Wgt_reg_279;
reg [18:0] Wgt_reg_280;
reg [18:0] Wgt_reg_281;
reg [18:0] Wgt_reg_282;
reg [18:0] Wgt_reg_283;
reg [18:0] Wgt_reg_284;
reg [18:0] Wgt_reg_285;
reg [18:0] Wgt_reg_286;
reg [18:0] Wgt_reg_287;
reg [18:0] Wgt_reg_288;
reg [18:0] Wgt_reg_289;
reg [18:0] Wgt_reg_290;
reg [18:0] Wgt_reg_291;
reg [18:0] Wgt_reg_292;
reg [18:0] Wgt_reg_293;
reg [18:0] Wgt_reg_294;
reg [18:0] Wgt_reg_295;
reg [18:0] Wgt_reg_296;
reg [18:0] Wgt_reg_297;
reg [18:0] Wgt_reg_298;
reg [18:0] Wgt_reg_299;
reg [18:0] Wgt_reg_300;
reg [18:0] Wgt_reg_301;
reg [18:0] Wgt_reg_302;
reg [18:0] Wgt_reg_303;
reg [18:0] Wgt_reg_304;
reg [18:0] Wgt_reg_305;
reg [18:0] Wgt_reg_306;
reg [18:0] Wgt_reg_307;
reg [18:0] Wgt_reg_308;
reg [18:0] Wgt_reg_309;
reg [18:0] Wgt_reg_310;
reg [18:0] Wgt_reg_311;
reg [18:0] Wgt_reg_312;
reg [18:0] Wgt_reg_313;
reg [18:0] Wgt_reg_314;
reg [18:0] Wgt_reg_315;
reg [18:0] Wgt_reg_316;
reg [18:0] Wgt_reg_317;
reg [18:0] Wgt_reg_318;
reg [18:0] Wgt_reg_319;
reg [18:0] Wgt_reg_320;
reg [18:0] Wgt_reg_321;
reg [18:0] Wgt_reg_322;
reg [18:0] Wgt_reg_323;
reg [18:0] Wgt_reg_324;
reg [18:0] Wgt_reg_325;
reg [18:0] Wgt_reg_326;
reg [18:0] Wgt_reg_327;
reg [18:0] Wgt_reg_328;
reg [18:0] Wgt_reg_329;
reg [18:0] Wgt_reg_330;
reg [18:0] Wgt_reg_331;
reg [18:0] Wgt_reg_332;
reg [18:0] Wgt_reg_333;
reg [18:0] Wgt_reg_334;
reg [18:0] Wgt_reg_335;
reg [18:0] Wgt_reg_336;
reg [18:0] Wgt_reg_337;
reg [18:0] Wgt_reg_338;
reg [18:0] Wgt_reg_339;
reg [18:0] Wgt_reg_340;
reg [18:0] Wgt_reg_341;
reg [18:0] Wgt_reg_342;
reg [18:0] Wgt_reg_343;
reg [18:0] Wgt_reg_344;
reg [18:0] Wgt_reg_345;
reg [18:0] Wgt_reg_346;
reg [18:0] Wgt_reg_347;
reg [18:0] Wgt_reg_348;
reg [18:0] Wgt_reg_349;
reg [18:0] Wgt_reg_350;
reg [18:0] Wgt_reg_351;
reg [18:0] Wgt_reg_352;
reg [18:0] Wgt_reg_353;
reg [18:0] Wgt_reg_354;
reg [18:0] Wgt_reg_355;
reg [18:0] Wgt_reg_356;
reg [18:0] Wgt_reg_357;
reg [18:0] Wgt_reg_358;
reg [18:0] Wgt_reg_359;
reg [18:0] Wgt_reg_360;
reg [18:0] Wgt_reg_361;
reg [18:0] Wgt_reg_362;
reg [18:0] Wgt_reg_363;
reg [18:0] Wgt_reg_364;
reg [18:0] Wgt_reg_365;
reg [18:0] Wgt_reg_366;
reg [18:0] Wgt_reg_367;
reg [18:0] Wgt_reg_368;
reg [18:0] Wgt_reg_369;
reg [18:0] Wgt_reg_370;
reg [18:0] Wgt_reg_371;
reg [18:0] Wgt_reg_372;
reg [18:0] Wgt_reg_373;
reg [18:0] Wgt_reg_374;
reg [18:0] Wgt_reg_375;
reg [18:0] Wgt_reg_376;
reg [18:0] Wgt_reg_377;
reg [18:0] Wgt_reg_378;
reg [18:0] Wgt_reg_379;
reg [18:0] Wgt_reg_380;
reg [18:0] Wgt_reg_381;
reg [18:0] Wgt_reg_382;
reg [18:0] Wgt_reg_383;
reg [18:0] Wgt_reg_384;
reg [18:0] Wgt_reg_385;
reg [18:0] Wgt_reg_386;
reg [18:0] Wgt_reg_387;
reg [18:0] Wgt_reg_388;
reg [18:0] Wgt_reg_389;
reg [18:0] Wgt_reg_390;
reg [18:0] Wgt_reg_391;
reg [18:0] Wgt_reg_392;
reg [18:0] Wgt_reg_393;
reg [18:0] Wgt_reg_394;
reg [18:0] Wgt_reg_395;
reg [18:0] Wgt_reg_396;
reg [18:0] Wgt_reg_397;
reg [18:0] Wgt_reg_398;
reg [18:0] Wgt_reg_399;
reg [18:0] Wgt_reg_400;
reg [18:0] Wgt_reg_401;
reg [18:0] Wgt_reg_402;
reg [18:0] Wgt_reg_403;
reg [18:0] Wgt_reg_404;
reg [18:0] Wgt_reg_405;
reg [18:0] Wgt_reg_406;
reg [18:0] Wgt_reg_407;
reg [18:0] Wgt_reg_408;
reg [18:0] Wgt_reg_409;
reg [18:0] Wgt_reg_410;
reg [18:0] Wgt_reg_411;
reg [18:0] Wgt_reg_412;
reg [18:0] Wgt_reg_413;
reg [18:0] Wgt_reg_414;
reg [18:0] Wgt_reg_415;
reg [18:0] Wgt_reg_416;
reg [18:0] Wgt_reg_417;
reg [18:0] Wgt_reg_418;
reg [18:0] Wgt_reg_419;
reg [18:0] Wgt_reg_420;
reg [18:0] Wgt_reg_421;
reg [18:0] Wgt_reg_422;
reg [18:0] Wgt_reg_423;
reg [18:0] Wgt_reg_424;
reg [18:0] Wgt_reg_425;
reg [18:0] Wgt_reg_426;
reg [18:0] Wgt_reg_427;
reg [18:0] Wgt_reg_428;
reg [18:0] Wgt_reg_429;
reg [18:0] Wgt_reg_430;
reg [18:0] Wgt_reg_431;
reg [18:0] Wgt_reg_432;
reg [18:0] Wgt_reg_433;
reg [18:0] Wgt_reg_434;
reg [18:0] Wgt_reg_435;
reg [18:0] Wgt_reg_436;
reg [18:0] Wgt_reg_437;
reg [18:0] Wgt_reg_438;
reg [18:0] Wgt_reg_439;
reg [18:0] Wgt_reg_440;
reg [18:0] Wgt_reg_441;
reg [18:0] Wgt_reg_442;
reg [18:0] Wgt_reg_443;
reg [18:0] Wgt_reg_444;
reg [18:0] Wgt_reg_445;
reg [18:0] Wgt_reg_446;
reg [18:0] Wgt_reg_447;
reg [18:0] Wgt_reg_448;
reg [18:0] Wgt_reg_449;
reg [18:0] Wgt_reg_450;
reg [18:0] Wgt_reg_451;
reg [18:0] Wgt_reg_452;
reg [18:0] Wgt_reg_453;
reg [18:0] Wgt_reg_454;
reg [18:0] Wgt_reg_455;
reg [18:0] Wgt_reg_456;
reg [18:0] Wgt_reg_457;
reg [18:0] Wgt_reg_458;
reg [18:0] Wgt_reg_459;
reg [18:0] Wgt_reg_460;
reg [18:0] Wgt_reg_461;
reg [18:0] Wgt_reg_462;
reg [18:0] Wgt_reg_463;
reg [18:0] Wgt_reg_464;
reg [18:0] Wgt_reg_465;
reg [18:0] Wgt_reg_466;
reg [18:0] Wgt_reg_467;
reg [18:0] Wgt_reg_468;
reg [18:0] Wgt_reg_469;
reg [18:0] Wgt_reg_470;
reg [18:0] Wgt_reg_471;
reg [18:0] Wgt_reg_472;
reg [18:0] Wgt_reg_473;
reg [18:0] Wgt_reg_474;
reg [18:0] Wgt_reg_475;
reg [18:0] Wgt_reg_476;
reg [18:0] Wgt_reg_477;
reg [18:0] Wgt_reg_478;
reg [18:0] Wgt_reg_479;
reg [18:0] Wgt_reg_480;
reg [18:0] Wgt_reg_481;
reg [18:0] Wgt_reg_482;
reg [18:0] Wgt_reg_483;
reg [18:0] Wgt_reg_484;
reg [18:0] Wgt_reg_485;
reg [18:0] Wgt_reg_486;
reg [18:0] Wgt_reg_487;
reg [18:0] Wgt_reg_488;
reg [18:0] Wgt_reg_489;
reg [18:0] Wgt_reg_490;
reg [18:0] Wgt_reg_491;
reg [18:0] Wgt_reg_492;
reg [18:0] Wgt_reg_493;
reg [18:0] Wgt_reg_494;
reg [18:0] Wgt_reg_495;
reg [18:0] Wgt_reg_496;
reg [18:0] Wgt_reg_497;
reg [18:0] Wgt_reg_498;
reg [18:0] Wgt_reg_499;
reg [18:0] Wgt_reg_500;
reg [18:0] Wgt_reg_501;
reg [18:0] Wgt_reg_502;
reg [18:0] Wgt_reg_503;
reg [18:0] Wgt_reg_504;
reg [18:0] Wgt_reg_505;
reg [18:0] Wgt_reg_506;
reg [18:0] Wgt_reg_507;
reg [18:0] Wgt_reg_508;
reg [18:0] Wgt_reg_509;
reg [18:0] Wgt_reg_510;
reg [18:0] Wgt_reg_511;
reg [18:0] Wgt_reg_512;
reg [18:0] Wgt_reg_513;
reg [18:0] Wgt_reg_514;
reg [18:0] Wgt_reg_515;
reg [18:0] Wgt_reg_516;
reg [18:0] Wgt_reg_517;
reg [18:0] Wgt_reg_518;
reg [18:0] Wgt_reg_519;
reg [18:0] Wgt_reg_520;
reg [18:0] Wgt_reg_521;
reg [18:0] Wgt_reg_522;
reg [18:0] Wgt_reg_523;
reg [18:0] Wgt_reg_524;
reg [18:0] Wgt_reg_525;
reg [18:0] Wgt_reg_526;
reg [18:0] Wgt_reg_527;
reg [18:0] Wgt_reg_528;
reg [18:0] Wgt_reg_529;
reg [18:0] Wgt_reg_530;
reg [18:0] Wgt_reg_531;
reg [18:0] Wgt_reg_532;
reg [18:0] Wgt_reg_533;
reg [18:0] Wgt_reg_534;
reg [18:0] Wgt_reg_535;
reg [18:0] Wgt_reg_536;
reg [18:0] Wgt_reg_537;
reg [18:0] Wgt_reg_538;
reg [18:0] Wgt_reg_539;
reg [18:0] Wgt_reg_540;
reg [18:0] Wgt_reg_541;
reg [18:0] Wgt_reg_542;
reg [18:0] Wgt_reg_543;
reg [18:0] Wgt_reg_544;
reg [18:0] Wgt_reg_545;
reg [18:0] Wgt_reg_546;
reg [18:0] Wgt_reg_547;
reg [18:0] Wgt_reg_548;
reg [18:0] Wgt_reg_549;
reg [18:0] Wgt_reg_550;
reg [18:0] Wgt_reg_551;
reg [18:0] Wgt_reg_552;
reg [18:0] Wgt_reg_553;
reg [18:0] Wgt_reg_554;
reg [18:0] Wgt_reg_555;
reg [18:0] Wgt_reg_556;
reg [18:0] Wgt_reg_557;
reg [18:0] Wgt_reg_558;
reg [18:0] Wgt_reg_559;
reg [18:0] Wgt_reg_560;
reg [18:0] Wgt_reg_561;
reg [18:0] Wgt_reg_562;
reg [18:0] Wgt_reg_563;
reg [18:0] Wgt_reg_564;
reg [18:0] Wgt_reg_565;
reg [18:0] Wgt_reg_566;
reg [18:0] Wgt_reg_567;
reg [18:0] Wgt_reg_568;
reg [18:0] Wgt_reg_569;
reg [18:0] Wgt_reg_570;
reg [18:0] Wgt_reg_571;
reg [18:0] Wgt_reg_572;
reg [18:0] Wgt_reg_573;
reg [18:0] Wgt_reg_574;
reg [18:0] Wgt_reg_575;
reg [18:0] Wgt_reg_576;
reg [18:0] Wgt_reg_577;
reg [18:0] Wgt_reg_578;
reg [18:0] Wgt_reg_579;
reg [18:0] Wgt_reg_580;
reg [18:0] Wgt_reg_581;
reg [18:0] Wgt_reg_582;
reg [18:0] Wgt_reg_583;
reg [18:0] Wgt_reg_584;
reg [18:0] Wgt_reg_585;
reg [18:0] Wgt_reg_586;
reg [18:0] Wgt_reg_587;
reg [18:0] Wgt_reg_588;
reg [18:0] Wgt_reg_589;
reg [18:0] Wgt_reg_590;
reg [18:0] Wgt_reg_591;
reg [18:0] Wgt_reg_592;
reg [18:0] Wgt_reg_593;
reg [18:0] Wgt_reg_594;
reg [18:0] Wgt_reg_595;
reg [18:0] Wgt_reg_596;
reg [18:0] Wgt_reg_597;
reg [18:0] Wgt_reg_598;
reg [18:0] Wgt_reg_599;
reg [18:0] Wgt_reg_600;
reg [18:0] Wgt_reg_601;
reg [18:0] Wgt_reg_602;
reg [18:0] Wgt_reg_603;
reg [18:0] Wgt_reg_604;
reg [18:0] Wgt_reg_605;
reg [18:0] Wgt_reg_606;
reg [18:0] Wgt_reg_607;
reg [18:0] Wgt_reg_608;
reg [18:0] Wgt_reg_609;
reg [18:0] Wgt_reg_610;
reg [18:0] Wgt_reg_611;
reg [18:0] Wgt_reg_612;
reg [18:0] Wgt_reg_613;
reg [18:0] Wgt_reg_614;
reg [18:0] Wgt_reg_615;
reg [18:0] Wgt_reg_616;
reg [18:0] Wgt_reg_617;
reg [18:0] Wgt_reg_618;
reg [18:0] Wgt_reg_619;
reg [18:0] Wgt_reg_620;
reg [18:0] Wgt_reg_621;
reg [18:0] Wgt_reg_622;
reg [18:0] Wgt_reg_623;
reg [18:0] Wgt_reg_624;
reg [18:0] Wgt_reg_625;
reg [18:0] Wgt_reg_626;
reg [18:0] Wgt_reg_627;
reg [18:0] Wgt_reg_628;
reg [18:0] Wgt_reg_629;
reg [18:0] Wgt_reg_630;
reg [18:0] Wgt_reg_631;
reg [18:0] Wgt_reg_632;
reg [18:0] Wgt_reg_633;
reg [18:0] Wgt_reg_634;
reg [18:0] Wgt_reg_635;
reg [18:0] Wgt_reg_636;
reg [18:0] Wgt_reg_637;
reg [18:0] Wgt_reg_638;
reg [18:0] Wgt_reg_639;
reg [18:0] Wgt_reg_640;
reg [18:0] Wgt_reg_641;
reg [18:0] Wgt_reg_642;
reg [18:0] Wgt_reg_643;
reg [18:0] Wgt_reg_644;
reg [18:0] Wgt_reg_645;
reg [18:0] Wgt_reg_646;
reg [18:0] Wgt_reg_647;
reg [18:0] Wgt_reg_648;
reg [18:0] Wgt_reg_649;
reg [18:0] Wgt_reg_650;
reg [18:0] Wgt_reg_651;
reg [18:0] Wgt_reg_652;
reg [18:0] Wgt_reg_653;
reg [18:0] Wgt_reg_654;
reg [18:0] Wgt_reg_655;
reg [18:0] Wgt_reg_656;
reg [18:0] Wgt_reg_657;
reg [18:0] Wgt_reg_658;
reg [18:0] Wgt_reg_659;
reg [18:0] Wgt_reg_660;
reg [18:0] Wgt_reg_661;
reg [18:0] Wgt_reg_662;
reg [18:0] Wgt_reg_663;
reg [18:0] Wgt_reg_664;
reg [18:0] Wgt_reg_665;
reg [18:0] Wgt_reg_666;
reg [18:0] Wgt_reg_667;
reg [18:0] Wgt_reg_668;
reg [18:0] Wgt_reg_669;
reg [18:0] Wgt_reg_670;
reg [18:0] Wgt_reg_671;
reg [18:0] Wgt_reg_672;
reg [18:0] Wgt_reg_673;
reg [18:0] Wgt_reg_674;
reg [18:0] Wgt_reg_675;
reg [18:0] Wgt_reg_676;
reg [18:0] Wgt_reg_677;
reg [18:0] Wgt_reg_678;
reg [18:0] Wgt_reg_679;
reg [18:0] Wgt_reg_680;
reg [18:0] Wgt_reg_681;
reg [18:0] Wgt_reg_682;
reg [18:0] Wgt_reg_683;
reg [18:0] Wgt_reg_684;
reg [18:0] Wgt_reg_685;
reg [18:0] Wgt_reg_686;
reg [18:0] Wgt_reg_687;
reg [18:0] Wgt_reg_688;
reg [18:0] Wgt_reg_689;
reg [18:0] Wgt_reg_690;
reg [18:0] Wgt_reg_691;
reg [18:0] Wgt_reg_692;
reg [18:0] Wgt_reg_693;
reg [18:0] Wgt_reg_694;
reg [18:0] Wgt_reg_695;
reg [18:0] Wgt_reg_696;
reg [18:0] Wgt_reg_697;
reg [18:0] Wgt_reg_698;
reg [18:0] Wgt_reg_699;
reg [18:0] Wgt_reg_700;
reg [18:0] Wgt_reg_701;
reg [18:0] Wgt_reg_702;
reg [18:0] Wgt_reg_703;
reg [18:0] Wgt_reg_704;
reg [18:0] Wgt_reg_705;
reg [18:0] Wgt_reg_706;
reg [18:0] Wgt_reg_707;
reg [18:0] Wgt_reg_708;
reg [18:0] Wgt_reg_709;
reg [18:0] Wgt_reg_710;
reg [18:0] Wgt_reg_711;
reg [18:0] Wgt_reg_712;
reg [18:0] Wgt_reg_713;
reg [18:0] Wgt_reg_714;
reg [18:0] Wgt_reg_715;
reg [18:0] Wgt_reg_716;
reg [18:0] Wgt_reg_717;
reg [18:0] Wgt_reg_718;
reg [18:0] Wgt_reg_719;
reg [18:0] Wgt_reg_720;
reg [18:0] Wgt_reg_721;
reg [18:0] Wgt_reg_722;
reg [18:0] Wgt_reg_723;
reg [18:0] Wgt_reg_724;
reg [18:0] Wgt_reg_725;
reg [18:0] Wgt_reg_726;
reg [18:0] Wgt_reg_727;
reg [18:0] Wgt_reg_728;
reg [18:0] Wgt_reg_729;
reg [18:0] Wgt_reg_730;
reg [18:0] Wgt_reg_731;
reg [18:0] Wgt_reg_732;
reg [18:0] Wgt_reg_733;
reg [18:0] Wgt_reg_734;
reg [18:0] Wgt_reg_735;
reg [18:0] Wgt_reg_736;
reg [18:0] Wgt_reg_737;
reg [18:0] Wgt_reg_738;
reg [18:0] Wgt_reg_739;
reg [18:0] Wgt_reg_740;
reg [18:0] Wgt_reg_741;
reg [18:0] Wgt_reg_742;
reg [18:0] Wgt_reg_743;
reg [18:0] Wgt_reg_744;
reg [18:0] Wgt_reg_745;
reg [18:0] Wgt_reg_746;
reg [18:0] Wgt_reg_747;
reg [18:0] Wgt_reg_748;
reg [18:0] Wgt_reg_749;
reg [18:0] Wgt_reg_750;
reg [18:0] Wgt_reg_751;
reg [18:0] Wgt_reg_752;
reg [18:0] Wgt_reg_753;
reg [18:0] Wgt_reg_754;
reg [18:0] Wgt_reg_755;
reg [18:0] Wgt_reg_756;
reg [18:0] Wgt_reg_757;
reg [18:0] Wgt_reg_758;
reg [18:0] Wgt_reg_759;
reg [18:0] Wgt_reg_760;
reg [18:0] Wgt_reg_761;
reg [18:0] Wgt_reg_762;
reg [18:0] Wgt_reg_763;
reg [18:0] Wgt_reg_764;
reg [18:0] Wgt_reg_765;
reg [18:0] Wgt_reg_766;
reg [18:0] Wgt_reg_767;
reg [18:0] Wgt_reg_768;
reg [18:0] Wgt_reg_769;
reg [18:0] Wgt_reg_770;
reg [18:0] Wgt_reg_771;
reg [18:0] Wgt_reg_772;
reg [18:0] Wgt_reg_773;
reg [18:0] Wgt_reg_774;
reg [18:0] Wgt_reg_775;
reg [18:0] Wgt_reg_776;
reg [18:0] Wgt_reg_777;
reg [18:0] Wgt_reg_778;
reg [18:0] Wgt_reg_779;
reg [18:0] Wgt_reg_780;
reg [18:0] Wgt_reg_781;
reg [18:0] Wgt_reg_782;
reg [18:0] Wgt_reg_783;
reg [18:0] Wgt_reg_784;




//mux pixels output  改成9位
wire [9:0] pixmuxout0;
wire [9:0] pixmuxout1;
wire [9:0] pixmuxout2;
wire [9:0] pixmuxout3;
wire [9:0] pixmuxout4;
wire [9:0] pixmuxout5;
wire [9:0] pixmuxout6;
wire [9:0] pixmuxout7;
wire [9:0] pixmuxout8;
wire [9:0] pixmuxout9;
wire [9:0] pixmuxout10;
wire [9:0] pixmuxout11;
wire [9:0] pixmuxout12;
wire [9:0] pixmuxout13;
wire [9:0] pixmuxout14;
wire [9:0] pixmuxout15;
wire [9:0] pixmuxout16;
wire [9:0] pixmuxout17;
wire [9:0] pixmuxout18;
wire [9:0] pixmuxout19;
wire [9:0] pixmuxout20;
wire [9:0] pixmuxout21;
wire [9:0] pixmuxout22;
wire [9:0] pixmuxout23;
wire [9:0] pixmuxout24;
wire [9:0] pixmuxout25;
wire [9:0] pixmuxout26;
wire [9:0] pixmuxout27;
//weight mux outputs 
wire [18:0] wtmuxout0;
wire [18:0] wtmuxout1;
wire [18:0] wtmuxout2;
wire [18:0] wtmuxout3;
wire [18:0] wtmuxout4;
wire [18:0] wtmuxout5;
wire [18:0] wtmuxout6;
wire [18:0] wtmuxout7;
wire [18:0] wtmuxout8;
wire [18:0] wtmuxout9;
wire [18:0] wtmuxout10;
wire [18:0] wtmuxout11;
wire [18:0] wtmuxout12;
wire [18:0] wtmuxout13;
wire [18:0] wtmuxout14;
wire [18:0] wtmuxout15;
wire [18:0] wtmuxout16;
wire [18:0] wtmuxout17;
wire [18:0] wtmuxout18;
wire [18:0] wtmuxout19;
wire [18:0] wtmuxout20;
wire [18:0] wtmuxout21;
wire [18:0] wtmuxout22;
wire [18:0] wtmuxout23;
wire [18:0] wtmuxout24;
wire [18:0] wtmuxout25;
wire [18:0] wtmuxout26;
wire [18:0] wtmuxout27;

//multiplier outputs
wire [25:0] multiout0;
wire [25:0] multiout1;
wire [25:0] multiout2;
wire [25:0] multiout3;
wire [25:0] multiout4;
wire [25:0] multiout5;
wire [25:0] multiout6;
wire [25:0] multiout7;
wire [25:0] multiout8;
wire [25:0] multiout9;
wire [25:0] multiout10;
wire [25:0] multiout11;
wire [25:0] multiout12;
wire [25:0] multiout13;
wire [25:0] multiout14;
wire [25:0] multiout15;
wire [25:0] multiout16;
wire [25:0] multiout17;
wire [25:0] multiout18;
wire [25:0] multiout19;
wire [25:0] multiout20;
wire [25:0] multiout21;
wire [25:0] multiout22;
wire [25:0] multiout23;
wire [25:0] multiout24;
wire [25:0] multiout25;
wire [25:0] multiout26;
wire [25:0] multiout27;

//1st level 14 adders' outputs
wire [25:0] addout0;
wire [25:0] addout1;
wire [25:0] addout2;
wire [25:0] addout3;
wire [25:0] addout4;
wire [25:0] addout5;
wire [25:0] addout6;
wire [25:0] addout7;
wire [25:0] addout8;
wire [25:0] addout9;
wire [25:0] addout10;
wire [25:0] addout11;
wire [25:0] addout12;
wire [25:0] addout13;

//2nd level 7 adders' outputs

wire [25:0] addout2nd_0;
wire [25:0] addout2nd_1;
wire [25:0] addout2nd_2;
wire [25:0] addout2nd_3;
wire [25:0] addout2nd_4;
wire [25:0] addout2nd_5;
wire [25:0] addout2nd_6;

//3rd level 4 adders' outputs (+ one more output from 2nd level passes the reg rather than adder)

wire [25:0] addout3rd_0;
wire [25:0] addout3rd_1;
wire [25:0] addout3rd_2;
wire [25:0] addout3rd_3;
//4th
wire [25:0] addout4th_0;
wire [25:0] addout4th_1;
//5th
wire [25:0] addout5th_0;
//total sum

wire [25:0] sum;

//bias
wire [25:0] bias;

//add all the sums
reg [25:0] zero_reg;
//1st level 14 add_sum_sumers' outputs
wire [25:0] add_sumout0;
wire [25:0] add_sumout1;
wire [25:0] add_sumout2;
wire [25:0] add_sumout3;
wire [25:0] add_sumout4;
wire [25:0] add_sumout5;
wire [25:0] add_sumout6;
wire [25:0] add_sumout7;
wire [25:0] add_sumout8;
wire [25:0] add_sumout9;
wire [25:0] add_sumout10;
wire [25:0] add_sumout11;
wire [25:0] add_sumout12;
wire [25:0] add_sumout13;

//2nd level 7 add_sumers' outputs

wire [25:0] add_sumout2nd_0;
wire [25:0] add_sumout2nd_1;
wire [25:0] add_sumout2nd_2;
wire [25:0] add_sumout2nd_3;
wire [25:0] add_sumout2nd_4;
wire [25:0] add_sumout2nd_5;
wire [25:0] add_sumout2nd_6;

//3rd level 4 add_sumers' outputs (+ one more output from 2nd level passes the reg rather than add_sumer)

wire [25:0] add_sumout3rd_0;
wire [25:0] add_sumout3rd_1;
wire [25:0] add_sumout3rd_2;
wire [25:0] add_sumout3rd_3;
//4th
wire [25:0] add_sumout4th_0;
wire [25:0] add_sumout4th_1;


muxpix mux0( //28to1 mux for pixels //可能还要加一个globalreset
select,
Pix_reg_0,
Pix_reg_1,
Pix_reg_2,
Pix_reg_3,
Pix_reg_4,
Pix_reg_5,
Pix_reg_6,
Pix_reg_7,
Pix_reg_8,
Pix_reg_9,
Pix_reg_10,
Pix_reg_11,
Pix_reg_12,
Pix_reg_13,
Pix_reg_14,
Pix_reg_15,
Pix_reg_16,
Pix_reg_17,
Pix_reg_18,
Pix_reg_19,
Pix_reg_20,
Pix_reg_21,
Pix_reg_22,
Pix_reg_23,
Pix_reg_24,
Pix_reg_25,
Pix_reg_26,
Pix_reg_27,
clk,
pixmuxout0
);

muxpix mux1( //28to1 mux for 
select,
Pix_reg_28,
Pix_reg_29,
Pix_reg_30,
Pix_reg_31,
Pix_reg_32,
Pix_reg_33,
Pix_reg_34,
Pix_reg_35,
Pix_reg_36,
Pix_reg_37,
Pix_reg_38,
Pix_reg_39,
Pix_reg_40,
Pix_reg_41,
Pix_reg_42,
Pix_reg_43,
Pix_reg_44,
Pix_reg_45,
Pix_reg_46,
Pix_reg_47,
Pix_reg_48,
Pix_reg_49,
Pix_reg_50,
Pix_reg_51,
Pix_reg_52,
Pix_reg_53,
Pix_reg_54,
Pix_reg_55,
clk,
pixmuxout1
);

muxpix mux2( //28to1 mux for 
select,
Pix_reg_56,
Pix_reg_57,
Pix_reg_58,
Pix_reg_59,
Pix_reg_60,
Pix_reg_61,
Pix_reg_62,
Pix_reg_63,
Pix_reg_64,
Pix_reg_65,
Pix_reg_66,
Pix_reg_67,
Pix_reg_68,
Pix_reg_69,
Pix_reg_70,
Pix_reg_71,
Pix_reg_72,
Pix_reg_73,
Pix_reg_74,
Pix_reg_75,
Pix_reg_76,
Pix_reg_77,
Pix_reg_78,
Pix_reg_79,
Pix_reg_80,
Pix_reg_81,
Pix_reg_82,
Pix_reg_83,
clk,
pixmuxout2
);

muxpix mux3( //28to1 mux for 
select,
Pix_reg_84,
Pix_reg_85,
Pix_reg_86,
Pix_reg_87,
Pix_reg_88,
Pix_reg_89,
Pix_reg_90,
Pix_reg_91,
Pix_reg_92,
Pix_reg_93,
Pix_reg_94,
Pix_reg_95,
Pix_reg_96,
Pix_reg_97,
Pix_reg_98,
Pix_reg_99,
Pix_reg_100,
Pix_reg_101,
Pix_reg_102,
Pix_reg_103,
Pix_reg_104,
Pix_reg_105,
Pix_reg_106,
Pix_reg_107,
Pix_reg_108,
Pix_reg_109,
Pix_reg_110,
Pix_reg_111,
clk,
pixmuxout3
);

muxpix mux4( //28to1 mux for weights
select,
Pix_reg_112,
Pix_reg_113,
Pix_reg_114,
Pix_reg_115,
Pix_reg_116,
Pix_reg_117,
Pix_reg_118,
Pix_reg_119,
Pix_reg_120,
Pix_reg_121,
Pix_reg_122,
Pix_reg_123,
Pix_reg_124,
Pix_reg_125,
Pix_reg_126,
Pix_reg_127,
Pix_reg_128,
Pix_reg_129,
Pix_reg_130,
Pix_reg_131,
Pix_reg_132,
Pix_reg_133,
Pix_reg_134,
Pix_reg_135,
Pix_reg_136,
Pix_reg_137,
Pix_reg_138,
Pix_reg_139,
clk,
pixmuxout4
);

muxpix mux5( //28to1 mux for weights
select,
Pix_reg_140,
Pix_reg_141,
Pix_reg_142,
Pix_reg_143,
Pix_reg_144,
Pix_reg_145,
Pix_reg_146,
Pix_reg_147,
Pix_reg_148,
Pix_reg_149,
Pix_reg_150,
Pix_reg_151,
Pix_reg_152,
Pix_reg_153,
Pix_reg_154,
Pix_reg_155,
Pix_reg_156,
Pix_reg_157,
Pix_reg_158,
Pix_reg_159,
Pix_reg_160,
Pix_reg_161,
Pix_reg_162,
Pix_reg_163,
Pix_reg_164,
Pix_reg_165,
Pix_reg_166,
Pix_reg_167,
clk,
pixmuxout5
);

muxpix mux6( //28to1 mux for weights
select,
Pix_reg_168,
Pix_reg_169,
Pix_reg_170,
Pix_reg_171,
Pix_reg_172,
Pix_reg_173,
Pix_reg_174,
Pix_reg_175,
Pix_reg_176,
Pix_reg_177,
Pix_reg_178,
Pix_reg_179,
Pix_reg_180,
Pix_reg_181,
Pix_reg_182,
Pix_reg_183,
Pix_reg_184,
Pix_reg_185,
Pix_reg_186,
Pix_reg_187,
Pix_reg_188,
Pix_reg_189,
Pix_reg_190,
Pix_reg_191,
Pix_reg_192,
Pix_reg_193,
Pix_reg_194,
Pix_reg_195,
clk,
pixmuxout6
);

muxpix mux7( //28to1 mux for weights
select,
Pix_reg_196,
Pix_reg_197,
Pix_reg_198,
Pix_reg_199,
Pix_reg_200,
Pix_reg_201,
Pix_reg_202,
Pix_reg_203,
Pix_reg_204,
Pix_reg_205,
Pix_reg_206,
Pix_reg_207,
Pix_reg_208,
Pix_reg_209,
Pix_reg_210,
Pix_reg_211,
Pix_reg_212,
Pix_reg_213,
Pix_reg_214,
Pix_reg_215,
Pix_reg_216,
Pix_reg_217,
Pix_reg_218,
Pix_reg_219,
Pix_reg_220,
Pix_reg_221,
Pix_reg_222,
Pix_reg_223,
clk,
pixmuxout7
);

muxpix mux8( //28to1 mux for weights
select,
Pix_reg_224,
Pix_reg_225,
Pix_reg_226,
Pix_reg_227,
Pix_reg_228,
Pix_reg_229,
Pix_reg_230,
Pix_reg_231,
Pix_reg_232,
Pix_reg_233,
Pix_reg_234,
Pix_reg_235,
Pix_reg_236,
Pix_reg_237,
Pix_reg_238,
Pix_reg_239,
Pix_reg_240,
Pix_reg_241,
Pix_reg_242,
Pix_reg_243,
Pix_reg_244,
Pix_reg_245,
Pix_reg_246,
Pix_reg_247,
Pix_reg_248,
Pix_reg_249,
Pix_reg_250,
Pix_reg_251,
clk,
pixmuxout8
);

muxpix mux9( //28to1 mux for weights
select,
Pix_reg_252,
Pix_reg_253,
Pix_reg_254,
Pix_reg_255,
Pix_reg_256,
Pix_reg_257,
Pix_reg_258,
Pix_reg_259,
Pix_reg_260,
Pix_reg_261,
Pix_reg_262,
Pix_reg_263,
Pix_reg_264,
Pix_reg_265,
Pix_reg_266,
Pix_reg_267,
Pix_reg_268,
Pix_reg_269,
Pix_reg_270,
Pix_reg_271,
Pix_reg_272,
Pix_reg_273,
Pix_reg_274,
Pix_reg_275,
Pix_reg_276,
Pix_reg_277,
Pix_reg_278,
Pix_reg_279,
clk,
pixmuxout9
);

muxpix mux10( //28to1 mux for weights
select,
Pix_reg_280,
Pix_reg_281,
Pix_reg_282,
Pix_reg_283,
Pix_reg_284,
Pix_reg_285,
Pix_reg_286,
Pix_reg_287,
Pix_reg_288,
Pix_reg_289,
Pix_reg_290,
Pix_reg_291,
Pix_reg_292,
Pix_reg_293,
Pix_reg_294,
Pix_reg_295,
Pix_reg_296,
Pix_reg_297,
Pix_reg_298,
Pix_reg_299,
Pix_reg_300,
Pix_reg_301,
Pix_reg_302,
Pix_reg_303,
Pix_reg_304,
Pix_reg_305,
Pix_reg_306,
Pix_reg_307,
clk,
pixmuxout10
);
muxpix mux11( //28to1 mux for weights
select,
Pix_reg_308,
Pix_reg_309,
Pix_reg_310,
Pix_reg_311,
Pix_reg_312,
Pix_reg_313,
Pix_reg_314,
Pix_reg_315,
Pix_reg_316,
Pix_reg_317,
Pix_reg_318,
Pix_reg_319,
Pix_reg_320,
Pix_reg_321,
Pix_reg_322,
Pix_reg_323,
Pix_reg_324,
Pix_reg_325,
Pix_reg_326,
Pix_reg_327,
Pix_reg_328,
Pix_reg_329,
Pix_reg_330,
Pix_reg_331,
Pix_reg_332,
Pix_reg_333,
Pix_reg_334,
Pix_reg_335,
clk,
pixmuxout11
);

muxpix mux12( //28to1 mux for weights
select,
Pix_reg_336,
Pix_reg_337,
Pix_reg_338,
Pix_reg_339,
Pix_reg_340,
Pix_reg_341,
Pix_reg_342,
Pix_reg_343,
Pix_reg_344,
Pix_reg_345,
Pix_reg_346,
Pix_reg_347,
Pix_reg_348,
Pix_reg_349,
Pix_reg_350,
Pix_reg_351,
Pix_reg_352,
Pix_reg_353,
Pix_reg_354,
Pix_reg_355,
Pix_reg_356,
Pix_reg_357,
Pix_reg_358,
Pix_reg_359,
Pix_reg_360,
Pix_reg_361,
Pix_reg_362,
Pix_reg_363,
clk,
pixmuxout12
);

muxpix mux13( //28to1 mux for weights
select,
Pix_reg_364,
Pix_reg_365,
Pix_reg_366,
Pix_reg_367,
Pix_reg_368,
Pix_reg_369,
Pix_reg_370,
Pix_reg_371,
Pix_reg_372,
Pix_reg_373,
Pix_reg_374,
Pix_reg_375,
Pix_reg_376,
Pix_reg_377,
Pix_reg_378,
Pix_reg_379,
Pix_reg_380,
Pix_reg_381,
Pix_reg_382,
Pix_reg_383,
Pix_reg_384,
Pix_reg_385,
Pix_reg_386,
Pix_reg_387,
Pix_reg_388,
Pix_reg_389,
Pix_reg_390,
Pix_reg_391,
clk,
pixmuxout13
);

muxpix mux14( //28to1 mux for weights
select,
Pix_reg_392,
Pix_reg_393,
Pix_reg_394,
Pix_reg_395,
Pix_reg_396,
Pix_reg_397,
Pix_reg_398,
Pix_reg_399,
Pix_reg_400,
Pix_reg_401,
Pix_reg_402,
Pix_reg_403,
Pix_reg_404,
Pix_reg_405,
Pix_reg_406,
Pix_reg_407,
Pix_reg_408,
Pix_reg_409,
Pix_reg_410,
Pix_reg_411,
Pix_reg_412,
Pix_reg_413,
Pix_reg_414,
Pix_reg_415,
Pix_reg_416,
Pix_reg_417,
Pix_reg_418,
Pix_reg_419,
clk,
pixmuxout14
);

muxpix mux15( //28to1 mux for weights
select,
Pix_reg_420,
Pix_reg_421,
Pix_reg_422,
Pix_reg_423,
Pix_reg_424,
Pix_reg_425,
Pix_reg_426,
Pix_reg_427,
Pix_reg_428,
Pix_reg_429,
Pix_reg_430,
Pix_reg_431,
Pix_reg_432,
Pix_reg_433,
Pix_reg_434,
Pix_reg_435,
Pix_reg_436,
Pix_reg_437,
Pix_reg_438,
Pix_reg_439,
Pix_reg_440,
Pix_reg_441,
Pix_reg_442,
Pix_reg_443,
Pix_reg_444,
Pix_reg_445,
Pix_reg_446,
Pix_reg_447,
clk,
pixmuxout15
);

muxpix mux16( //28to1 mux for weights
select,
Pix_reg_448,
Pix_reg_449,
Pix_reg_450,
Pix_reg_451,
Pix_reg_452,
Pix_reg_453,
Pix_reg_454,
Pix_reg_455,
Pix_reg_456,
Pix_reg_457,
Pix_reg_458,
Pix_reg_459,
Pix_reg_460,
Pix_reg_461,
Pix_reg_462,
Pix_reg_463,
Pix_reg_464,
Pix_reg_465,
Pix_reg_466,
Pix_reg_467,
Pix_reg_468,
Pix_reg_469,
Pix_reg_470,
Pix_reg_471,
Pix_reg_472,
Pix_reg_473,
Pix_reg_474,
Pix_reg_475,
clk,
pixmuxout16
);

muxpix mux17( //28to1 mux for weights
select,
Pix_reg_476,
Pix_reg_477,
Pix_reg_478,
Pix_reg_479,
Pix_reg_480,
Pix_reg_481,
Pix_reg_482,
Pix_reg_483,
Pix_reg_484,
Pix_reg_485,
Pix_reg_486,
Pix_reg_487,
Pix_reg_488,
Pix_reg_489,
Pix_reg_490,
Pix_reg_491,
Pix_reg_492,
Pix_reg_493,
Pix_reg_494,
Pix_reg_495,
Pix_reg_496,
Pix_reg_497,
Pix_reg_498,
Pix_reg_499,
Pix_reg_500,
Pix_reg_501,
Pix_reg_502,
Pix_reg_503,
clk,
pixmuxout17
);

muxpix mux18( //28to1 mux for weights
select,
Pix_reg_504,
Pix_reg_505,
Pix_reg_506,
Pix_reg_507,
Pix_reg_508,
Pix_reg_509,
Pix_reg_510,
Pix_reg_511,
Pix_reg_512,
Pix_reg_513,
Pix_reg_514,
Pix_reg_515,
Pix_reg_516,
Pix_reg_517,
Pix_reg_518,
Pix_reg_519,
Pix_reg_520,
Pix_reg_521,
Pix_reg_522,
Pix_reg_523,
Pix_reg_524,
Pix_reg_525,
Pix_reg_526,
Pix_reg_527,
Pix_reg_528,
Pix_reg_529,
Pix_reg_530,
Pix_reg_531,
clk,
pixmuxout18
);

muxpix mux19( //28to1 mux for weights
select,
Pix_reg_532,
Pix_reg_533,
Pix_reg_534,
Pix_reg_535,
Pix_reg_536,
Pix_reg_537,
Pix_reg_538,
Pix_reg_539,
Pix_reg_540,
Pix_reg_541,
Pix_reg_542,
Pix_reg_543,
Pix_reg_544,
Pix_reg_545,
Pix_reg_546,
Pix_reg_547,
Pix_reg_548,
Pix_reg_549,
Pix_reg_550,
Pix_reg_551,
Pix_reg_552,
Pix_reg_553,
Pix_reg_554,
Pix_reg_555,
Pix_reg_556,
Pix_reg_557,
Pix_reg_558,
Pix_reg_559,
clk,
pixmuxout19
);

muxpix mux20( //28to1 mux for weights
select,
Pix_reg_560,
Pix_reg_561,
Pix_reg_562,
Pix_reg_563,
Pix_reg_564,
Pix_reg_565,
Pix_reg_566,
Pix_reg_567,
Pix_reg_568,
Pix_reg_569,
Pix_reg_570,
Pix_reg_571,
Pix_reg_572,
Pix_reg_573,
Pix_reg_574,
Pix_reg_575,
Pix_reg_576,
Pix_reg_577,
Pix_reg_578,
Pix_reg_579,
Pix_reg_580,
Pix_reg_581,
Pix_reg_582,
Pix_reg_583,
Pix_reg_584,
Pix_reg_585,
Pix_reg_586,
Pix_reg_587,
clk,
pixmuxout20
);
muxpix mux21( //28to1 mux for weights
select,
Pix_reg_588,
Pix_reg_589,
Pix_reg_590,
Pix_reg_591,
Pix_reg_592,
Pix_reg_593,
Pix_reg_594,
Pix_reg_595,
Pix_reg_596,
Pix_reg_597,
Pix_reg_598,
Pix_reg_599,
Pix_reg_600,
Pix_reg_601,
Pix_reg_602,
Pix_reg_603,
Pix_reg_604,
Pix_reg_605,
Pix_reg_606,
Pix_reg_607,
Pix_reg_608,
Pix_reg_609,
Pix_reg_610,
Pix_reg_611,
Pix_reg_612,
Pix_reg_613,
Pix_reg_614,
Pix_reg_615,
clk,
pixmuxout21
);

muxpix mux22( //28to1 mux for weights
select,
Pix_reg_616,
Pix_reg_617,
Pix_reg_618,
Pix_reg_619,
Pix_reg_620,
Pix_reg_621,
Pix_reg_622,
Pix_reg_623,
Pix_reg_624,
Pix_reg_625,
Pix_reg_626,
Pix_reg_627,
Pix_reg_628,
Pix_reg_629,
Pix_reg_630,
Pix_reg_631,
Pix_reg_632,
Pix_reg_633,
Pix_reg_634,
Pix_reg_635,
Pix_reg_636,
Pix_reg_637,
Pix_reg_638,
Pix_reg_639,
Pix_reg_640,
Pix_reg_641,
Pix_reg_642,
Pix_reg_643,
clk,
pixmuxout22
);

muxpix mux23( //28to1 mux for weights
select,
Pix_reg_644,
Pix_reg_645,
Pix_reg_646,
Pix_reg_647,
Pix_reg_648,
Pix_reg_649,
Pix_reg_650,
Pix_reg_651,
Pix_reg_652,
Pix_reg_653,
Pix_reg_654,
Pix_reg_655,
Pix_reg_656,
Pix_reg_657,
Pix_reg_658,
Pix_reg_659,
Pix_reg_660,
Pix_reg_661,
Pix_reg_662,
Pix_reg_663,
Pix_reg_664,
Pix_reg_665,
Pix_reg_666,
Pix_reg_667,
Pix_reg_668,
Pix_reg_669,
Pix_reg_670,
Pix_reg_671,
clk,
pixmuxout23
);

muxpix mux24( //28to1 mux for weights
select,
Pix_reg_672,
Pix_reg_673,
Pix_reg_674,
Pix_reg_675,
Pix_reg_676,
Pix_reg_677,
Pix_reg_678,
Pix_reg_679,
Pix_reg_680,
Pix_reg_681,
Pix_reg_682,
Pix_reg_683,
Pix_reg_684,
Pix_reg_685,
Pix_reg_686,
Pix_reg_687,
Pix_reg_688,
Pix_reg_689,
Pix_reg_690,
Pix_reg_691,
Pix_reg_692,
Pix_reg_693,
Pix_reg_694,
Pix_reg_695,
Pix_reg_696,
Pix_reg_697,
Pix_reg_698,
Pix_reg_699,
clk,
pixmuxout24
);

muxpix mux25( //28to1 mux for weights
select,
Pix_reg_700,
Pix_reg_701,
Pix_reg_702,
Pix_reg_703,
Pix_reg_704,
Pix_reg_705,
Pix_reg_706,
Pix_reg_707,
Pix_reg_708,
Pix_reg_709,
Pix_reg_710,
Pix_reg_711,
Pix_reg_712,
Pix_reg_713,
Pix_reg_714,
Pix_reg_715,
Pix_reg_716,
Pix_reg_717,
Pix_reg_718,
Pix_reg_719,
Pix_reg_720,
Pix_reg_721,
Pix_reg_722,
Pix_reg_723,
Pix_reg_724,
Pix_reg_725,
Pix_reg_726,
Pix_reg_727,
clk,
pixmuxout25
);
muxpix mux26( //28to1 mux for weights
select,
Pix_reg_728,
Pix_reg_729,
Pix_reg_730,
Pix_reg_731,
Pix_reg_732,
Pix_reg_733,
Pix_reg_734,
Pix_reg_735,
Pix_reg_736,
Pix_reg_737,
Pix_reg_738,
Pix_reg_739,
Pix_reg_740,
Pix_reg_741,
Pix_reg_742,
Pix_reg_743,
Pix_reg_744,
Pix_reg_745,
Pix_reg_746,
Pix_reg_747,
Pix_reg_748,
Pix_reg_749,
Pix_reg_750,
Pix_reg_751,
Pix_reg_752,
Pix_reg_753,
Pix_reg_754,
Pix_reg_755,
clk,
pixmuxout26
);

muxpix mux27( //28to1 mux for weights
select,
Pix_reg_756,
Pix_reg_757,
Pix_reg_758,
Pix_reg_759,
Pix_reg_760,
Pix_reg_761,
Pix_reg_762,
Pix_reg_763,
Pix_reg_764,
Pix_reg_765,
Pix_reg_766,
Pix_reg_767,
Pix_reg_768,
Pix_reg_769,
Pix_reg_770,
Pix_reg_771,
Pix_reg_772,
Pix_reg_773,
Pix_reg_774,
Pix_reg_775,
Pix_reg_776,
Pix_reg_777,
Pix_reg_778,
Pix_reg_779,
Pix_reg_780,
Pix_reg_781,
Pix_reg_782,
Pix_reg_783,
clk,
pixmuxout27
);


mux wtmux0( //28to1 mux for  
select,
 Wgt_reg_0,
 Wgt_reg_1,
 Wgt_reg_2,
 Wgt_reg_3,
 Wgt_reg_4,
 Wgt_reg_5,
 Wgt_reg_6,
 Wgt_reg_7,
 Wgt_reg_8,
 Wgt_reg_9,
 Wgt_reg_10,
 Wgt_reg_11,
 Wgt_reg_12,
 Wgt_reg_13,
 Wgt_reg_14,
 Wgt_reg_15,
 Wgt_reg_16,
 Wgt_reg_17,
 Wgt_reg_18,
 Wgt_reg_19,
 Wgt_reg_20,
 Wgt_reg_21,
 Wgt_reg_22,
 Wgt_reg_23,
 Wgt_reg_24,
 Wgt_reg_25,
 Wgt_reg_26,
 Wgt_reg_27,
clk,
wtmuxout0
);

mux wtmux1( //28to1 mux for 
 select,
 Wgt_reg_28,
 Wgt_reg_29,
 Wgt_reg_30,
 Wgt_reg_31,
 Wgt_reg_32,
 Wgt_reg_33,
 Wgt_reg_34,
 Wgt_reg_35,
 Wgt_reg_36,
 Wgt_reg_37,
 Wgt_reg_38,
 Wgt_reg_39,
 Wgt_reg_40,
 Wgt_reg_41,
 Wgt_reg_42,
 Wgt_reg_43,
 Wgt_reg_44,
 Wgt_reg_45,
 Wgt_reg_46,
 Wgt_reg_47,
 Wgt_reg_48,
 Wgt_reg_49,
 Wgt_reg_50,
 Wgt_reg_51,
 Wgt_reg_52,
 Wgt_reg_53,
 Wgt_reg_54,
 Wgt_reg_55,
clk,
wtmuxout1
);

mux wtmux2( //28to1 mux for 
select,
 Wgt_reg_56,
 Wgt_reg_57,
 Wgt_reg_58,
 Wgt_reg_59,
 Wgt_reg_60,
 Wgt_reg_61,
 Wgt_reg_62,
 Wgt_reg_63,
 Wgt_reg_64,
 Wgt_reg_65,
 Wgt_reg_66,
 Wgt_reg_67,
 Wgt_reg_68,
 Wgt_reg_69,
 Wgt_reg_70,
 Wgt_reg_71,
 Wgt_reg_72,
 Wgt_reg_73,
 Wgt_reg_74,
 Wgt_reg_75,
 Wgt_reg_76,
 Wgt_reg_77,
 Wgt_reg_78,
 Wgt_reg_79,
 Wgt_reg_80,
 Wgt_reg_81,
 Wgt_reg_82,
 Wgt_reg_83,
clk,
wtmuxout2
);

mux wtmux3( //28to1 mux for 
select,
 Wgt_reg_84,
 Wgt_reg_85,
 Wgt_reg_86,
 Wgt_reg_87,
 Wgt_reg_88,
 Wgt_reg_89,
 Wgt_reg_90,
 Wgt_reg_91,
 Wgt_reg_92,
 Wgt_reg_93,
 Wgt_reg_94,
 Wgt_reg_95,
 Wgt_reg_96,
 Wgt_reg_97,
 Wgt_reg_98,
 Wgt_reg_99,
 Wgt_reg_100,
 Wgt_reg_101,
 Wgt_reg_102,
 Wgt_reg_103,
 Wgt_reg_104,
 Wgt_reg_105,
 Wgt_reg_106,
 Wgt_reg_107,
 Wgt_reg_108,
 Wgt_reg_109,
 Wgt_reg_110,
 Wgt_reg_111,
clk,
wtmuxout3
);

mux wtmux4( //28to1 mux for weights
select,
 Wgt_reg_112,
 Wgt_reg_113,
 Wgt_reg_114,
 Wgt_reg_115,
 Wgt_reg_116,
 Wgt_reg_117,
 Wgt_reg_118,
 Wgt_reg_119,
 Wgt_reg_120,
 Wgt_reg_121,
 Wgt_reg_122,
 Wgt_reg_123,
 Wgt_reg_124,
 Wgt_reg_125,
 Wgt_reg_126,
 Wgt_reg_127,
 Wgt_reg_128,
 Wgt_reg_129,
 Wgt_reg_130,
 Wgt_reg_131,
 Wgt_reg_132,
 Wgt_reg_133,
 Wgt_reg_134,
 Wgt_reg_135,
 Wgt_reg_136,
 Wgt_reg_137,
 Wgt_reg_138,
 Wgt_reg_139,
clk,
wtmuxout4
);

mux wtmux5( //28to1 mux for weights
select,
 Wgt_reg_140,
 Wgt_reg_141,
 Wgt_reg_142,
 Wgt_reg_143,
 Wgt_reg_144,
 Wgt_reg_145,
 Wgt_reg_146,
 Wgt_reg_147,
 Wgt_reg_148,
 Wgt_reg_149,
 Wgt_reg_150,
 Wgt_reg_151,
 Wgt_reg_152,
 Wgt_reg_153,
 Wgt_reg_154,
 Wgt_reg_155,
 Wgt_reg_156,
 Wgt_reg_157,
 Wgt_reg_158,
 Wgt_reg_159,
 Wgt_reg_160,
 Wgt_reg_161,
 Wgt_reg_162,
 Wgt_reg_163,
 Wgt_reg_164,
 Wgt_reg_165,
 Wgt_reg_166,
 Wgt_reg_167,
clk,
wtmuxout5
);

mux wtmux6( //28to1 mux for weights
select,
 Wgt_reg_168,
 Wgt_reg_169,
 Wgt_reg_170,
 Wgt_reg_171,
 Wgt_reg_172,
 Wgt_reg_173,
 Wgt_reg_174,
 Wgt_reg_175,
 Wgt_reg_176,
 Wgt_reg_177,
 Wgt_reg_178,
 Wgt_reg_179,
 Wgt_reg_180,
 Wgt_reg_181,
 Wgt_reg_182,
 Wgt_reg_183,
 Wgt_reg_184,
 Wgt_reg_185,
 Wgt_reg_186,
 Wgt_reg_187,
 Wgt_reg_188,
 Wgt_reg_189,
 Wgt_reg_190,
 Wgt_reg_191,
 Wgt_reg_192,
 Wgt_reg_193,
 Wgt_reg_194,
 Wgt_reg_195,
clk,
wtmuxout6
);

mux wtmux7( //28to1 mux for weights
select,
 Wgt_reg_196,
 Wgt_reg_197,
 Wgt_reg_198,
 Wgt_reg_199,
 Wgt_reg_200,
 Wgt_reg_201,
 Wgt_reg_202,
 Wgt_reg_203,
 Wgt_reg_204,
 Wgt_reg_205,
 Wgt_reg_206,
 Wgt_reg_207,
 Wgt_reg_208,
 Wgt_reg_209,
 Wgt_reg_210,
 Wgt_reg_211,
 Wgt_reg_212,
 Wgt_reg_213,
 Wgt_reg_214,
 Wgt_reg_215,
 Wgt_reg_216,
 Wgt_reg_217,
 Wgt_reg_218,
 Wgt_reg_219,
 Wgt_reg_220,
 Wgt_reg_221,
 Wgt_reg_222,
 Wgt_reg_223,
clk,
wtmuxout7
);

mux wtmux8( //28to1 mux for weights
select,
 Wgt_reg_224,
 Wgt_reg_225,
 Wgt_reg_226,
 Wgt_reg_227,
 Wgt_reg_228,
 Wgt_reg_229,
 Wgt_reg_230,
 Wgt_reg_231,
 Wgt_reg_232,
 Wgt_reg_233,
 Wgt_reg_234,
 Wgt_reg_235,
 Wgt_reg_236,
 Wgt_reg_237,
 Wgt_reg_238,
 Wgt_reg_239,
 Wgt_reg_240,
 Wgt_reg_241,
 Wgt_reg_242,
 Wgt_reg_243,
 Wgt_reg_244,
 Wgt_reg_245,
 Wgt_reg_246,
 Wgt_reg_247,
 Wgt_reg_248,
 Wgt_reg_249,
 Wgt_reg_250,
 Wgt_reg_251,
clk,
wtmuxout8
);

mux wtmux9( //28to1 mux for weights
select,
 Wgt_reg_252,
 Wgt_reg_253,
 Wgt_reg_254,
 Wgt_reg_255,
 Wgt_reg_256,
 Wgt_reg_257,
 Wgt_reg_258,
 Wgt_reg_259,
 Wgt_reg_260,
 Wgt_reg_261,
 Wgt_reg_262,
 Wgt_reg_263,
 Wgt_reg_264,
 Wgt_reg_265,
 Wgt_reg_266,
 Wgt_reg_267,
 Wgt_reg_268,
 Wgt_reg_269,
 Wgt_reg_270,
 Wgt_reg_271,
 Wgt_reg_272,
 Wgt_reg_273,
 Wgt_reg_274,
 Wgt_reg_275,
 Wgt_reg_276,
 Wgt_reg_277,
 Wgt_reg_278,
 Wgt_reg_279,
clk,
wtmuxout9
);

mux wtmux10( //28to1 mux for weights
select,
 Wgt_reg_280,
 Wgt_reg_281,
 Wgt_reg_282,
 Wgt_reg_283,
 Wgt_reg_284,
 Wgt_reg_285,
 Wgt_reg_286,
 Wgt_reg_287,
 Wgt_reg_288,
 Wgt_reg_289,
 Wgt_reg_290,
 Wgt_reg_291,
 Wgt_reg_292,
 Wgt_reg_293,
 Wgt_reg_294,
 Wgt_reg_295,
 Wgt_reg_296,
 Wgt_reg_297,
 Wgt_reg_298,
 Wgt_reg_299,
 Wgt_reg_300,
 Wgt_reg_301,
 Wgt_reg_302,
 Wgt_reg_303,
 Wgt_reg_304,
 Wgt_reg_305,
 Wgt_reg_306,
 Wgt_reg_307,
clk,
wtmuxout10
);
mux wtmux11( //28to1 mux for weights
select,
 Wgt_reg_308,
 Wgt_reg_309,
 Wgt_reg_310,
 Wgt_reg_311,
 Wgt_reg_312,
 Wgt_reg_313,
 Wgt_reg_314,
 Wgt_reg_315,
 Wgt_reg_316,
 Wgt_reg_317,
 Wgt_reg_318,
 Wgt_reg_319,
 Wgt_reg_320,
 Wgt_reg_321,
 Wgt_reg_322,
 Wgt_reg_323,
 Wgt_reg_324,
 Wgt_reg_325,
 Wgt_reg_326,
 Wgt_reg_327,
 Wgt_reg_328,
 Wgt_reg_329,
 Wgt_reg_330,
 Wgt_reg_331,
 Wgt_reg_332,
 Wgt_reg_333,
 Wgt_reg_334,
 Wgt_reg_335,
clk,
wtmuxout11
);

mux wtmux12( //28to1 mux for weights
select,
 Wgt_reg_336,
 Wgt_reg_337,
 Wgt_reg_338,
 Wgt_reg_339,
 Wgt_reg_340,
 Wgt_reg_341,
 Wgt_reg_342,
 Wgt_reg_343,
 Wgt_reg_344,
 Wgt_reg_345,
 Wgt_reg_346,
 Wgt_reg_347,
 Wgt_reg_348,
 Wgt_reg_349,
 Wgt_reg_350,
 Wgt_reg_351,
 Wgt_reg_352,
 Wgt_reg_353,
 Wgt_reg_354,
 Wgt_reg_355,
 Wgt_reg_356,
 Wgt_reg_357,
 Wgt_reg_358,
 Wgt_reg_359,
 Wgt_reg_360,
 Wgt_reg_361,
 Wgt_reg_362,
 Wgt_reg_363,
clk,
wtmuxout12
);

mux wtmux13( //28to1 mux for weights
select,
 Wgt_reg_364,
 Wgt_reg_365,
 Wgt_reg_366,
 Wgt_reg_367,
 Wgt_reg_368,
 Wgt_reg_369,
 Wgt_reg_370,
 Wgt_reg_371,
 Wgt_reg_372,
 Wgt_reg_373,
 Wgt_reg_374,
 Wgt_reg_375,
 Wgt_reg_376,
 Wgt_reg_377,
 Wgt_reg_378,
 Wgt_reg_379,
 Wgt_reg_380,
 Wgt_reg_381,
 Wgt_reg_382,
 Wgt_reg_383,
 Wgt_reg_384,
 Wgt_reg_385,
 Wgt_reg_386,
 Wgt_reg_387,
 Wgt_reg_388,
 Wgt_reg_389,
 Wgt_reg_390,
 Wgt_reg_391,
clk,
wtmuxout13
);

mux wtmux14( //28to1 mux for weights
select,
 Wgt_reg_392,
 Wgt_reg_393,
 Wgt_reg_394,
 Wgt_reg_395,
 Wgt_reg_396,
 Wgt_reg_397,
 Wgt_reg_398,
 Wgt_reg_399,
 Wgt_reg_400,
 Wgt_reg_401,
 Wgt_reg_402,
 Wgt_reg_403,
 Wgt_reg_404,
 Wgt_reg_405,
 Wgt_reg_406,
 Wgt_reg_407,
 Wgt_reg_408,
 Wgt_reg_409,
 Wgt_reg_410,
 Wgt_reg_411,
 Wgt_reg_412,
 Wgt_reg_413,
 Wgt_reg_414,
 Wgt_reg_415,
 Wgt_reg_416,
 Wgt_reg_417,
 Wgt_reg_418,
 Wgt_reg_419,
clk,
wtmuxout14
);

mux wtmux15( //28to1 mux for weights
select,
 Wgt_reg_420,
 Wgt_reg_421,
 Wgt_reg_422,
 Wgt_reg_423,
 Wgt_reg_424,
 Wgt_reg_425,
 Wgt_reg_426,
 Wgt_reg_427,
 Wgt_reg_428,
 Wgt_reg_429,
 Wgt_reg_430,
 Wgt_reg_431,
 Wgt_reg_432,
 Wgt_reg_433,
 Wgt_reg_434,
 Wgt_reg_435,
 Wgt_reg_436,
 Wgt_reg_437,
 Wgt_reg_438,
 Wgt_reg_439,
 Wgt_reg_440,
 Wgt_reg_441,
 Wgt_reg_442,
 Wgt_reg_443,
 Wgt_reg_444,
 Wgt_reg_445,
 Wgt_reg_446,
 Wgt_reg_447,
clk,
wtmuxout15
);

mux wtmux16( //28to1 mux for weights
select,
 Wgt_reg_448,
 Wgt_reg_449,
 Wgt_reg_450,
 Wgt_reg_451,
 Wgt_reg_452,
 Wgt_reg_453,
 Wgt_reg_454,
 Wgt_reg_455,
 Wgt_reg_456,
 Wgt_reg_457,
 Wgt_reg_458,
 Wgt_reg_459,
 Wgt_reg_460,
 Wgt_reg_461,
 Wgt_reg_462,
 Wgt_reg_463,
 Wgt_reg_464,
 Wgt_reg_465,
 Wgt_reg_466,
 Wgt_reg_467,
 Wgt_reg_468,
 Wgt_reg_469,
 Wgt_reg_470,
 Wgt_reg_471,
 Wgt_reg_472,
 Wgt_reg_473,
 Wgt_reg_474,
 Wgt_reg_475,
clk,
wtmuxout16
);

mux wtmux17( //28to1 mux for weights
select,
 Wgt_reg_476,
 Wgt_reg_477,
 Wgt_reg_478,
 Wgt_reg_479,
 Wgt_reg_480,
 Wgt_reg_481,
 Wgt_reg_482,
 Wgt_reg_483,
 Wgt_reg_484,
 Wgt_reg_485,
 Wgt_reg_486,
 Wgt_reg_487,
 Wgt_reg_488,
 Wgt_reg_489,
 Wgt_reg_490,
 Wgt_reg_491,
 Wgt_reg_492,
 Wgt_reg_493,
 Wgt_reg_494,
 Wgt_reg_495,
 Wgt_reg_496,
 Wgt_reg_497,
 Wgt_reg_498,
 Wgt_reg_499,
 Wgt_reg_500,
 Wgt_reg_501,
 Wgt_reg_502,
 Wgt_reg_503,
clk,
wtmuxout17
);

mux wtmux18( //28to1 mux for weights
select,
 Wgt_reg_504,
 Wgt_reg_505,
 Wgt_reg_506,
 Wgt_reg_507,
 Wgt_reg_508,
 Wgt_reg_509,
 Wgt_reg_510,
 Wgt_reg_511,
 Wgt_reg_512,
 Wgt_reg_513,
 Wgt_reg_514,
 Wgt_reg_515,
 Wgt_reg_516,
 Wgt_reg_517,
 Wgt_reg_518,
 Wgt_reg_519,
 Wgt_reg_520,
 Wgt_reg_521,
 Wgt_reg_522,
 Wgt_reg_523,
 Wgt_reg_524,
 Wgt_reg_525,
 Wgt_reg_526,
 Wgt_reg_527,
 Wgt_reg_528,
 Wgt_reg_529,
 Wgt_reg_530,
 Wgt_reg_531,
clk,
wtmuxout18
);

mux wtmux19( //28to1 mux for weights
select,
 Wgt_reg_532,
 Wgt_reg_533,
 Wgt_reg_534,
 Wgt_reg_535,
 Wgt_reg_536,
 Wgt_reg_537,
 Wgt_reg_538,
 Wgt_reg_539,
 Wgt_reg_540,
 Wgt_reg_541,
 Wgt_reg_542,
 Wgt_reg_543,
 Wgt_reg_544,
 Wgt_reg_545,
 Wgt_reg_546,
 Wgt_reg_547,
 Wgt_reg_548,
 Wgt_reg_549,
 Wgt_reg_550,
 Wgt_reg_551,
 Wgt_reg_552,
 Wgt_reg_553,
 Wgt_reg_554,
 Wgt_reg_555,
 Wgt_reg_556,
 Wgt_reg_557,
 Wgt_reg_558,
 Wgt_reg_559,
clk,
wtmuxout19
);

mux wtmux20( //28to1 mux for weights
select,
 Wgt_reg_560,
 Wgt_reg_561,
 Wgt_reg_562,
 Wgt_reg_563,
 Wgt_reg_564,
 Wgt_reg_565,
 Wgt_reg_566,
 Wgt_reg_567,
 Wgt_reg_568,
 Wgt_reg_569,
 Wgt_reg_570,
 Wgt_reg_571,
 Wgt_reg_572,
 Wgt_reg_573,
 Wgt_reg_574,
 Wgt_reg_575,
 Wgt_reg_576,
 Wgt_reg_577,
 Wgt_reg_578,
 Wgt_reg_579,
 Wgt_reg_580,
 Wgt_reg_581,
 Wgt_reg_582,
 Wgt_reg_583,
 Wgt_reg_584,
 Wgt_reg_585,
 Wgt_reg_586,
 Wgt_reg_587,
clk,
wtmuxout20
);
mux wtmux21( //28to1 mux for weights
select,
 Wgt_reg_588,
 Wgt_reg_589,
 Wgt_reg_590,
 Wgt_reg_591,
 Wgt_reg_592,
 Wgt_reg_593,
 Wgt_reg_594,
 Wgt_reg_595,
 Wgt_reg_596,
 Wgt_reg_597,
 Wgt_reg_598,
 Wgt_reg_599,
 Wgt_reg_600,
 Wgt_reg_601,
 Wgt_reg_602,
 Wgt_reg_603,
 Wgt_reg_604,
 Wgt_reg_605,
 Wgt_reg_606,
 Wgt_reg_607,
 Wgt_reg_608,
 Wgt_reg_609,
 Wgt_reg_610,
 Wgt_reg_611,
 Wgt_reg_612,
 Wgt_reg_613,
 Wgt_reg_614,
 Wgt_reg_615,
clk,
wtmuxout21
);

mux wtmux22( //28to1 mux for weights
select,
 Wgt_reg_616,
 Wgt_reg_617,
 Wgt_reg_618,
 Wgt_reg_619,
 Wgt_reg_620,
 Wgt_reg_621,
 Wgt_reg_622,
 Wgt_reg_623,
 Wgt_reg_624,
 Wgt_reg_625,
 Wgt_reg_626,
 Wgt_reg_627,
 Wgt_reg_628,
 Wgt_reg_629,
 Wgt_reg_630,
 Wgt_reg_631,
 Wgt_reg_632,
 Wgt_reg_633,
 Wgt_reg_634,
 Wgt_reg_635,
 Wgt_reg_636,
 Wgt_reg_637,
 Wgt_reg_638,
 Wgt_reg_639,
 Wgt_reg_640,
 Wgt_reg_641,
 Wgt_reg_642,
 Wgt_reg_643,
clk,
wtmuxout22
);

mux wtmux23( //28to1 mux for weights
select,
 Wgt_reg_644,
 Wgt_reg_645,
 Wgt_reg_646,
 Wgt_reg_647,
 Wgt_reg_648,
 Wgt_reg_649,
 Wgt_reg_650,
 Wgt_reg_651,
 Wgt_reg_652,
 Wgt_reg_653,
 Wgt_reg_654,
 Wgt_reg_655,
 Wgt_reg_656,
 Wgt_reg_657,
 Wgt_reg_658,
 Wgt_reg_659,
 Wgt_reg_660,
 Wgt_reg_661,
 Wgt_reg_662,
 Wgt_reg_663,
 Wgt_reg_664,
 Wgt_reg_665,
 Wgt_reg_666,
 Wgt_reg_667,
 Wgt_reg_668,
 Wgt_reg_669,
 Wgt_reg_670,
 Wgt_reg_671,
clk,
wtmuxout23
);

mux wtmux24( //28to1 mux for weights
select,
 Wgt_reg_672,
 Wgt_reg_673,
 Wgt_reg_674,
 Wgt_reg_675,
 Wgt_reg_676,
 Wgt_reg_677,
 Wgt_reg_678,
 Wgt_reg_679,
 Wgt_reg_680,
 Wgt_reg_681,
 Wgt_reg_682,
 Wgt_reg_683,
 Wgt_reg_684,
 Wgt_reg_685,
 Wgt_reg_686,
 Wgt_reg_687,
 Wgt_reg_688,
 Wgt_reg_689,
 Wgt_reg_690,
 Wgt_reg_691,
 Wgt_reg_692,
 Wgt_reg_693,
 Wgt_reg_694,
 Wgt_reg_695,
 Wgt_reg_696,
 Wgt_reg_697,
 Wgt_reg_698,
 Wgt_reg_699,
clk,
wtmuxout24
);

mux wtmux25( //28to1 mux for weights
select,
 Wgt_reg_700,
 Wgt_reg_701,
 Wgt_reg_702,
 Wgt_reg_703,
 Wgt_reg_704,
 Wgt_reg_705,
 Wgt_reg_706,
 Wgt_reg_707,
 Wgt_reg_708,
 Wgt_reg_709,
 Wgt_reg_710,
 Wgt_reg_711,
 Wgt_reg_712,
 Wgt_reg_713,
 Wgt_reg_714,
 Wgt_reg_715,
 Wgt_reg_716,
 Wgt_reg_717,
 Wgt_reg_718,
 Wgt_reg_719,
 Wgt_reg_720,
 Wgt_reg_721,
 Wgt_reg_722,
 Wgt_reg_723,
 Wgt_reg_724,
 Wgt_reg_725,
 Wgt_reg_726,
 Wgt_reg_727,
clk,
wtmuxout25
);
mux wtmux26( //28to1 mux for weights
select,
 Wgt_reg_728,
 Wgt_reg_729,
 Wgt_reg_730,
 Wgt_reg_731,
 Wgt_reg_732,
 Wgt_reg_733,
 Wgt_reg_734,
 Wgt_reg_735,
 Wgt_reg_736,
 Wgt_reg_737,
 Wgt_reg_738,
 Wgt_reg_739,
 Wgt_reg_740,
 Wgt_reg_741,
 Wgt_reg_742,
 Wgt_reg_743,
 Wgt_reg_744,
 Wgt_reg_745,
 Wgt_reg_746,
 Wgt_reg_747,
 Wgt_reg_748,
 Wgt_reg_749,
 Wgt_reg_750,
 Wgt_reg_751,
 Wgt_reg_752,
 Wgt_reg_753,
 Wgt_reg_754,
 Wgt_reg_755,
clk,
wtmuxout26
);

mux wtmux27( //28to1 mux for weights
select,
 Wgt_reg_756,
 Wgt_reg_757,
 Wgt_reg_758,
 Wgt_reg_759,
 Wgt_reg_760,
 Wgt_reg_761,
 Wgt_reg_762,
 Wgt_reg_763,
 Wgt_reg_764,
 Wgt_reg_765,
 Wgt_reg_766,
 Wgt_reg_767,
 Wgt_reg_768,
 Wgt_reg_769,
 Wgt_reg_770,
 Wgt_reg_771,
 Wgt_reg_772,
 Wgt_reg_773,
 Wgt_reg_774,
 Wgt_reg_775,
 Wgt_reg_776,
 Wgt_reg_777,
 Wgt_reg_778,
 Wgt_reg_779,
 Wgt_reg_780,
 Wgt_reg_781,
 Wgt_reg_782,
 Wgt_reg_783,
clk,
wtmuxout27
);

//mux for pixel还没写！！！
FixedPointMultiplier multi0 (
  clk,
  ~GlobalReset,
  wtmuxout0, // sfix19_En18
  pixmuxout0, // sfix10_En0
  multiout0 // sfix26_En18

);

FixedPointMultiplier multi1(
clk,
~GlobalReset,
 wtmuxout1,
pixmuxout1,
multiout1
	);

FixedPointMultiplier multi2(
clk,
~GlobalReset,
 wtmuxout2,
pixmuxout2,
multiout2
	);

FixedPointMultiplier multi3(
clk,
~GlobalReset,
 wtmuxout3,
pixmuxout3,
multiout3
	);

FixedPointMultiplier multi4(
clk,
~GlobalReset,
 wtmuxout4,
pixmuxout4,
multiout4
	);

FixedPointMultiplier multi5(
clk,
~GlobalReset,
 wtmuxout5,
pixmuxout5,
multiout5
	);

FixedPointMultiplier multi6(
clk,
~GlobalReset,
 wtmuxout6,
pixmuxout6,
multiout6
	);

FixedPointMultiplier multi7(
clk,
~GlobalReset,
 wtmuxout7,
pixmuxout7,
multiout7
	);

FixedPointMultiplier multi8(
clk,
~GlobalReset,
wtmuxout8,
pixmuxout8,
multiout8
	);

FixedPointMultiplier multi9(
clk,
~GlobalReset,
 wtmuxout9,
pixmuxout9,
multiout9
	);

FixedPointMultiplier multi10(
clk,
~GlobalReset,
 wtmuxout10,
pixmuxout10,
multiout10
	);

FixedPointMultiplier multi11(
clk,
~GlobalReset,
 wtmuxout11,
pixmuxout11,
multiout11
	);

FixedPointMultiplier multi12(
clk,
~GlobalReset,
 wtmuxout12,
pixmuxout12,
multiout12
	);

FixedPointMultiplier multi13(
clk,
~GlobalReset,
 wtmuxout13,
pixmuxout13,
multiout13
	);

FixedPointMultiplier multi14(
clk,
~GlobalReset,
 wtmuxout14,
pixmuxout14,
multiout14
	);

FixedPointMultiplier multi15(
clk,
~GlobalReset,
 wtmuxout15,
pixmuxout15,
multiout15
	);

FixedPointMultiplier multi16(
clk,
~GlobalReset,
 wtmuxout16,
pixmuxout16,
multiout16
	);

FixedPointMultiplier multi17(
clk,
~GlobalReset,
 wtmuxout17,
pixmuxout17,
multiout17
	);

FixedPointMultiplier multi18(
clk,
~GlobalReset,
 wtmuxout18,
pixmuxout18,
multiout18
	);

FixedPointMultiplier multi19(
clk,
~GlobalReset,
 wtmuxout19,
pixmuxout19,
multiout19
	);

FixedPointMultiplier multi20(
clk,
~GlobalReset,
 wtmuxout20,
pixmuxout20,
multiout20
	);

FixedPointMultiplier multi21(
clk,
~GlobalReset,
 wtmuxout21,
pixmuxout21,
multiout21
	);

FixedPointMultiplier multi22(
clk,
~GlobalReset,
 wtmuxout22,
pixmuxout22,
multiout22
	);

FixedPointMultiplier multi23(
clk,
~GlobalReset,
 wtmuxout23,
pixmuxout23,
multiout23
	);

FixedPointMultiplier multi24(
clk,
~GlobalReset,
 wtmuxout24,
pixmuxout24,
multiout24
	);

FixedPointMultiplier multi25(
clk,
~GlobalReset,
 wtmuxout25,
pixmuxout25,
multiout25
	);

FixedPointMultiplier multi26(
clk,
~GlobalReset,
 wtmuxout26,
pixmuxout26,
multiout26
);

FixedPointMultiplier multi27(
clk,
~GlobalReset,
 wtmuxout27,
pixmuxout27,
multiout27
);


FixedPointMultiplier multi_bias(
clk,
~GlobalReset,
Wgt_reg_784,
Pix_reg_784,
bias
);


FixedPointAdder add0(
  clk,
  ~GlobalReset,
  multiout0, 
  multiout1, 
  addout0
);

FixedPointAdder add1(
clk,
~GlobalReset,
multiout2, 
multiout3, 
addout1
	);

FixedPointAdder add2(
clk,
~GlobalReset,
multiout4, 
multiout5, 
addout2
	);

FixedPointAdder add3(
clk,
~GlobalReset,
multiout6, 
multiout7, 
addout3
	);

FixedPointAdder add4(
clk,
~GlobalReset,
multiout8, 
multiout9, 
addout4
	);

FixedPointAdder add5(
clk,
~GlobalReset,
multiout10, 
multiout11, 
addout5
	);

FixedPointAdder add6(
clk,
~GlobalReset,
multiout12, 
multiout13, 
addout6
	);

FixedPointAdder add7(
clk,
~GlobalReset,
multiout14, 
multiout15, 
addout7
	);

FixedPointAdder add8(
clk,
~GlobalReset,
multiout16, 
multiout17, 
addout8
	);

FixedPointAdder add9(
clk,
~GlobalReset,
multiout18, 
multiout19, 
addout9
	);

FixedPointAdder add10(
clk,
~GlobalReset,
multiout20, 
multiout21, 
addout10
	);

FixedPointAdder add11(
clk,
~GlobalReset,
multiout22, 
multiout23, 
addout11
	);

FixedPointAdder add12(
clk,
~GlobalReset,
multiout24, 
multiout25, 
addout12
	);

FixedPointAdder add13(
clk,
~GlobalReset,
multiout26, 
multiout27, 
addout13
	);


FixedPointAdder add2nd_0(
clk,
~GlobalReset,
addout0, 
addout1, 
addout2nd_0
	);

FixedPointAdder add2nd_1(
clk,
~GlobalReset,
addout2, 
addout3, 
addout2nd_1
	);

FixedPointAdder add2nd_2(
clk,
~GlobalReset,
addout4, 
addout5, 
addout2nd_2
	);

FixedPointAdder add2nd_3(
clk,
~GlobalReset,
addout6, 
addout7, 
addout2nd_3
	);

FixedPointAdder add2nd_4(
clk,
~GlobalReset,
addout8, 
addout9, 
addout2nd_4
	);

FixedPointAdder add2nd_5(
clk,
~GlobalReset,
addout10, 
addout11, 
addout2nd_5
	);

FixedPointAdder add2nd_6(
clk,
~GlobalReset,
addout12, 
addout13, 
addout2nd_6
	);

//addout3rd_0

FixedPointAdder add3rd_0(
clk,
~GlobalReset,
addout2nd_0, 
addout2nd_1, 
addout3rd_0
	);

FixedPointAdder add3rd_1(
clk,
~GlobalReset,
addout2nd_2, 
addout2nd_3, 
addout3rd_1
	);
FixedPointAdder add3rd_2(
clk,
~GlobalReset,
addout2nd_4, 
addout2nd_5, 
addout3rd_2
	);

FixedPointAdder add3rd_3(  //7th addout from 2nd level and the bias beta
clk,
~GlobalReset,
addout2nd_6, 
//{{(7){Wgt_784[18]}},Wgt_784},// or zero_reg, 
//{7'b0000000,Wgt_784},
//bias,
zero_reg,
addout3rd_3
	);


FixedPointAdder add4th_0(
clk,
~GlobalReset,
addout3rd_0, 
addout3rd_1, 
addout4th_0
	);

FixedPointAdder add4th_1(
clk,
~GlobalReset,
addout3rd_2, 
addout3rd_3, //
addout4th_1
	);

FixedPointAdder add5th_0(
clk,
~GlobalReset,
addout4th_0, 
addout4th_1, 
sum//addout5th_0
	);


FixedPointAdder add_sum0(
  clk,
  ~GlobalReset,
  sum_sim_reg0, 
  sum_sim_reg1, 
  add_sumout0
);

FixedPointAdder add_sum1(
clk,
~GlobalReset,
sum_sim_reg2, 
sum_sim_reg3, 
add_sumout1
	);

FixedPointAdder add_sum2(
clk,
~GlobalReset,
sum_sim_reg4, 
sum_sim_reg5, 
add_sumout2
	);

FixedPointAdder add_sum3(
clk,
~GlobalReset,
sum_sim_reg6, 
sum_sim_reg7, 
add_sumout3
	);

FixedPointAdder add_sum4(
clk,
~GlobalReset,
sum_sim_reg8, 
sum_sim_reg9, 
add_sumout4
	);

FixedPointAdder add_sum5(
clk,
~GlobalReset,
sum_sim_reg10, 
sum_sim_reg11, 
add_sumout5
	);

FixedPointAdder add_sum6(
clk,
~GlobalReset,
sum_sim_reg12, 
sum_sim_reg13, 
add_sumout6
	);

FixedPointAdder add_sum7(
clk,
~GlobalReset,
sum_sim_reg14, 
sum_sim_reg15, 
add_sumout7
	);

FixedPointAdder add_sum8(
clk,
~GlobalReset,
sum_sim_reg16, 
sum_sim_reg17, 
add_sumout8
	);

FixedPointAdder add_sum9(
clk,
~GlobalReset,
sum_sim_reg18, 
sum_sim_reg19, 
add_sumout9
	);

FixedPointAdder add_sum10(
clk,
~GlobalReset,
sum_sim_reg20, 
sum_sim_reg21, 
add_sumout10
	);

FixedPointAdder add_sum11(
clk,
~GlobalReset,
sum_sim_reg22, 
sum_sim_reg23, 
add_sumout11
	);

FixedPointAdder add_sum12(
clk,
~GlobalReset,
sum_sim_reg24, 
sum_sim_reg25, 
add_sumout12
	);

FixedPointAdder add_sum13(
clk,
~GlobalReset,
sum_sim_reg26, 
sum_sim_reg27, 
add_sumout13
	);


FixedPointAdder add_sum2nd_0(
clk,
~GlobalReset,
add_sumout0, 
add_sumout1, 
add_sumout2nd_0
	);

FixedPointAdder add_sum2nd_1(
clk,
~GlobalReset,
add_sumout2, 
add_sumout3, 
add_sumout2nd_1
	);

FixedPointAdder add_sum2nd_2(
clk,
~GlobalReset,
add_sumout4, 
add_sumout5, 
add_sumout2nd_2
	);

FixedPointAdder add_sum2nd_3(
clk,
~GlobalReset,
add_sumout6, 
add_sumout7, 
add_sumout2nd_3
	);

FixedPointAdder add_sum2nd_4(
clk,
~GlobalReset,
add_sumout8, 
add_sumout9, 
add_sumout2nd_4
	);

FixedPointAdder add_sum2nd_5(
clk,
~GlobalReset,
add_sumout10, 
add_sumout11, 
add_sumout2nd_5
	);

FixedPointAdder add_sum2nd_6(
clk,
~GlobalReset,
add_sumout12, 
add_sumout13, 
add_sumout2nd_6
	);

//add_sumout3rd_0

FixedPointAdder add_sum3rd_0(
clk,
~GlobalReset,
add_sumout2nd_0, 
add_sumout2nd_1, 
add_sumout3rd_0
	);

FixedPointAdder add_sum3rd_1(
clk,
~GlobalReset,
add_sumout2nd_2, 
add_sumout2nd_3, 
add_sumout3rd_1
	);
FixedPointAdder add_sum3rd_2(
clk,
~GlobalReset,
add_sumout2nd_4, 
add_sumout2nd_5, 
add_sumout3rd_2
	);

FixedPointAdder add_sum3rd_3(  //7th add_sumout from 2nd level and the bias beta
clk,
~GlobalReset,
add_sumout2nd_6, 
zero_reg,
add_sumout3rd_3
	);


FixedPointAdder add_sum4th_0(
clk,
~GlobalReset,
add_sumout3rd_0, 
add_sumout3rd_1, 
add_sumout4th_0
	);

FixedPointAdder add_sum4th_1(
clk,
~GlobalReset,
add_sumout3rd_2, 
add_sumout3rd_3, //
add_sumout4th_1
	);

FixedPointAdder add_sum5th_0(
clk,
~GlobalReset,
add_sumout4th_0, 
add_sumout4th_1, 
tot_out
	);

FixedPointAdder add_last(
clk,
~GlobalReset,
tot_out, 
bias,
tot_out_real
	);


/*FixedPointAdder addbias(
clk,
GlobalReset,
addout5th_0, 
Wgt_784, 
sum
	);*/
//reg[25:0] tot_out_r;
//assign tot_out = tot_out_r;

always @(posedge clk) begin 
	if (GlobalReset==0) begin
		state<=7'b0000000;
		
		
	end
	else begin
	case(state)
		7'b0000000: begin
		   Output_Valid_r<=1'b0;
		   if (Input_Valid==1)begin
			//select<=6'b000000;
			//Output_Valid_r <= 1'b0;
			zero_reg <= 26'b00000000000000000000000000;
			sum_sim_reg0 <=0;
         sum_sim_reg1 <=0;
         sum_sim_reg2 <=0;
         sum_sim_reg3 <=0;
         sum_sim_reg4 <=0;
         sum_sim_reg5 <=0;
         sum_sim_reg6 <=0;
         sum_sim_reg7 <=0;
         sum_sim_reg8 <=0;
         sum_sim_reg9 <=0;
         sum_sim_reg10 <=0;
         sum_sim_reg11 <=0;
         sum_sim_reg12 <=0;
      	 sum_sim_reg13 <=0;
         sum_sim_reg14 <=0;
         sum_sim_reg15 <=0;
         sum_sim_reg16 <=0;
         sum_sim_reg17 <=0;
         sum_sim_reg18 <=0;
         sum_sim_reg19 <=0;
         sum_sim_reg20 <=0;
         sum_sim_reg21 <=0;
         sum_sim_reg22 <=0;
         sum_sim_reg23 <=0;
         sum_sim_reg24 <=0;
         sum_sim_reg25 <=0;
         sum_sim_reg26 <=0;
         sum_sim_reg27 <=0;
		 cell_out_r<=0;


		Pix_reg_0 <= Pix_0;
		Pix_reg_1 <= Pix_1;
		Pix_reg_2 <= Pix_2;
		Pix_reg_3 <= Pix_3;
		Pix_reg_4 <= Pix_4;
		Pix_reg_5 <= Pix_5;
		Pix_reg_6 <= Pix_6;
		Pix_reg_7 <= Pix_7;
		Pix_reg_8 <= Pix_8;
		Pix_reg_9 <= Pix_9;
		Pix_reg_10 <= Pix_10;
		Pix_reg_11 <= Pix_11;
		Pix_reg_12 <= Pix_12;
		Pix_reg_13 <= Pix_13;
		Pix_reg_14 <= Pix_14;
		Pix_reg_15 <= Pix_15;
		Pix_reg_16 <= Pix_16;
		Pix_reg_17 <= Pix_17;
		Pix_reg_18 <= Pix_18;
		Pix_reg_19 <= Pix_19;
		Pix_reg_20 <= Pix_20;
		Pix_reg_21 <= Pix_21;
		Pix_reg_22 <= Pix_22;
		Pix_reg_23 <= Pix_23;
		Pix_reg_24 <= Pix_24;
		Pix_reg_25 <= Pix_25;
		Pix_reg_26 <= Pix_26;
		Pix_reg_27 <= Pix_27;
		Pix_reg_28 <= Pix_28;
		Pix_reg_29 <= Pix_29;
		Pix_reg_30 <= Pix_30;
		Pix_reg_31 <= Pix_31;
		Pix_reg_32 <= Pix_32;
		Pix_reg_33 <= Pix_33;
		Pix_reg_34 <= Pix_34;
		Pix_reg_35 <= Pix_35;
		Pix_reg_36 <= Pix_36;
		Pix_reg_37 <= Pix_37;
		Pix_reg_38 <= Pix_38;
		Pix_reg_39 <= Pix_39;
		Pix_reg_40 <= Pix_40;
		Pix_reg_41 <= Pix_41;
		Pix_reg_42 <= Pix_42;
		Pix_reg_43 <= Pix_43;
		Pix_reg_44 <= Pix_44;
		Pix_reg_45 <= Pix_45;
		Pix_reg_46 <= Pix_46;
		Pix_reg_47 <= Pix_47;
		Pix_reg_48 <= Pix_48;
		Pix_reg_49 <= Pix_49;
		Pix_reg_50 <= Pix_50;
		Pix_reg_51 <= Pix_51;
		Pix_reg_52 <= Pix_52;
		Pix_reg_53 <= Pix_53;
		Pix_reg_54 <= Pix_54;
		Pix_reg_55 <= Pix_55;
		Pix_reg_56 <= Pix_56;
		Pix_reg_57 <= Pix_57;
		Pix_reg_58 <= Pix_58;
		Pix_reg_59 <= Pix_59;
		Pix_reg_60 <= Pix_60;
		Pix_reg_61 <= Pix_61;
		Pix_reg_62 <= Pix_62;
		Pix_reg_63 <= Pix_63;
		Pix_reg_64 <= Pix_64;
		Pix_reg_65 <= Pix_65;
		Pix_reg_66 <= Pix_66;
		Pix_reg_67 <= Pix_67;
		Pix_reg_68 <= Pix_68;
		Pix_reg_69 <= Pix_69;
		Pix_reg_70 <= Pix_70;
		Pix_reg_71 <= Pix_71;
		Pix_reg_72 <= Pix_72;
		Pix_reg_73 <= Pix_73;
		Pix_reg_74 <= Pix_74;
		Pix_reg_75 <= Pix_75;
		Pix_reg_76 <= Pix_76;
		Pix_reg_77 <= Pix_77;
		Pix_reg_78 <= Pix_78;
		Pix_reg_79 <= Pix_79;
		Pix_reg_80 <= Pix_80;
		Pix_reg_81 <= Pix_81;
		Pix_reg_82 <= Pix_82;
		Pix_reg_83 <= Pix_83;
		Pix_reg_84 <= Pix_84;
		Pix_reg_85 <= Pix_85;
		Pix_reg_86 <= Pix_86;
		Pix_reg_87 <= Pix_87;
		Pix_reg_88 <= Pix_88;
		Pix_reg_89 <= Pix_89;
		Pix_reg_90 <= Pix_90;
		Pix_reg_91 <= Pix_91;
		Pix_reg_92 <= Pix_92;
		Pix_reg_93 <= Pix_93;
		Pix_reg_94 <= Pix_94;
		Pix_reg_95 <= Pix_95;
		Pix_reg_96 <= Pix_96;
		Pix_reg_97 <= Pix_97;
		Pix_reg_98 <= Pix_98;
		Pix_reg_99 <= Pix_99;
		Pix_reg_100 <= Pix_100;
		Pix_reg_101 <= Pix_101;
		Pix_reg_102 <= Pix_102;
		Pix_reg_103 <= Pix_103;
		Pix_reg_104 <= Pix_104;
		Pix_reg_105 <= Pix_105;
		Pix_reg_106 <= Pix_106;
		Pix_reg_107 <= Pix_107;
		Pix_reg_108 <= Pix_108;
		Pix_reg_109 <= Pix_109;
		Pix_reg_110 <= Pix_110;
		Pix_reg_111 <= Pix_111;
		Pix_reg_112 <= Pix_112;
		Pix_reg_113 <= Pix_113;
		Pix_reg_114 <= Pix_114;
		Pix_reg_115 <= Pix_115;
		Pix_reg_116 <= Pix_116;
		Pix_reg_117 <= Pix_117;
		Pix_reg_118 <= Pix_118;
		Pix_reg_119 <= Pix_119;
		Pix_reg_120 <= Pix_120;
		Pix_reg_121 <= Pix_121;
		Pix_reg_122 <= Pix_122;
		Pix_reg_123 <= Pix_123;
		Pix_reg_124 <= Pix_124;
		Pix_reg_125 <= Pix_125;
		Pix_reg_126 <= Pix_126;
		Pix_reg_127 <= Pix_127;
		Pix_reg_128 <= Pix_128;
		Pix_reg_129 <= Pix_129;
		Pix_reg_130 <= Pix_130;
		Pix_reg_131 <= Pix_131;
		Pix_reg_132 <= Pix_132;
		Pix_reg_133 <= Pix_133;
		Pix_reg_134 <= Pix_134;
		Pix_reg_135 <= Pix_135;
		Pix_reg_136 <= Pix_136;
		Pix_reg_137 <= Pix_137;
		Pix_reg_138 <= Pix_138;
		Pix_reg_139 <= Pix_139;
		Pix_reg_140 <= Pix_140;
		Pix_reg_141 <= Pix_141;
		Pix_reg_142 <= Pix_142;
		Pix_reg_143 <= Pix_143;
		Pix_reg_144 <= Pix_144;
		Pix_reg_145 <= Pix_145;
		Pix_reg_146 <= Pix_146;
		Pix_reg_147 <= Pix_147;
		Pix_reg_148 <= Pix_148;
		Pix_reg_149 <= Pix_149;
		Pix_reg_150 <= Pix_150;
		Pix_reg_151 <= Pix_151;
		Pix_reg_152 <= Pix_152;
		Pix_reg_153 <= Pix_153;
		Pix_reg_154 <= Pix_154;
		Pix_reg_155 <= Pix_155;
		Pix_reg_156 <= Pix_156;
		Pix_reg_157 <= Pix_157;
		Pix_reg_158 <= Pix_158;
		Pix_reg_159 <= Pix_159;
		Pix_reg_160 <= Pix_160;
		Pix_reg_161 <= Pix_161;
		Pix_reg_162 <= Pix_162;
		Pix_reg_163 <= Pix_163;
		Pix_reg_164 <= Pix_164;
		Pix_reg_165 <= Pix_165;
		Pix_reg_166 <= Pix_166;
		Pix_reg_167 <= Pix_167;
		Pix_reg_168 <= Pix_168;
		Pix_reg_169 <= Pix_169;
		Pix_reg_170 <= Pix_170;
		Pix_reg_171 <= Pix_171;
		Pix_reg_172 <= Pix_172;
		Pix_reg_173 <= Pix_173;
		Pix_reg_174 <= Pix_174;
		Pix_reg_175 <= Pix_175;
		Pix_reg_176 <= Pix_176;
		Pix_reg_177 <= Pix_177;
		Pix_reg_178 <= Pix_178;
		Pix_reg_179 <= Pix_179;
		Pix_reg_180 <= Pix_180;
		Pix_reg_181 <= Pix_181;
		Pix_reg_182 <= Pix_182;
		Pix_reg_183 <= Pix_183;
		Pix_reg_184 <= Pix_184;
		Pix_reg_185 <= Pix_185;
		Pix_reg_186 <= Pix_186;
		Pix_reg_187 <= Pix_187;
		Pix_reg_188 <= Pix_188;
		Pix_reg_189 <= Pix_189;
		Pix_reg_190 <= Pix_190;
		Pix_reg_191 <= Pix_191;
		Pix_reg_192 <= Pix_192;
		Pix_reg_193 <= Pix_193;
		Pix_reg_194 <= Pix_194;
		Pix_reg_195 <= Pix_195;
		Pix_reg_196 <= Pix_196;
		Pix_reg_197 <= Pix_197;
		Pix_reg_198 <= Pix_198;
		Pix_reg_199 <= Pix_199;
		Pix_reg_200 <= Pix_200;
		Pix_reg_201 <= Pix_201;
		Pix_reg_202 <= Pix_202;
		Pix_reg_203 <= Pix_203;
		Pix_reg_204 <= Pix_204;
		Pix_reg_205 <= Pix_205;
		Pix_reg_206 <= Pix_206;
		Pix_reg_207 <= Pix_207;
		Pix_reg_208 <= Pix_208;
		Pix_reg_209 <= Pix_209;
		Pix_reg_210 <= Pix_210;
		Pix_reg_211 <= Pix_211;
		Pix_reg_212 <= Pix_212;
		Pix_reg_213 <= Pix_213;
		Pix_reg_214 <= Pix_214;
		Pix_reg_215 <= Pix_215;
		Pix_reg_216 <= Pix_216;
		Pix_reg_217 <= Pix_217;
		Pix_reg_218 <= Pix_218;
		Pix_reg_219 <= Pix_219;
		Pix_reg_220 <= Pix_220;
		Pix_reg_221 <= Pix_221;
		Pix_reg_222 <= Pix_222;
		Pix_reg_223 <= Pix_223;
		Pix_reg_224 <= Pix_224;
		Pix_reg_225 <= Pix_225;
		Pix_reg_226 <= Pix_226;
		Pix_reg_227 <= Pix_227;
		Pix_reg_228 <= Pix_228;
		Pix_reg_229 <= Pix_229;
		Pix_reg_230 <= Pix_230;
		Pix_reg_231 <= Pix_231;
		Pix_reg_232 <= Pix_232;
		Pix_reg_233 <= Pix_233;
		Pix_reg_234 <= Pix_234;
		Pix_reg_235 <= Pix_235;
		Pix_reg_236 <= Pix_236;
		Pix_reg_237 <= Pix_237;
		Pix_reg_238 <= Pix_238;
		Pix_reg_239 <= Pix_239;
		Pix_reg_240 <= Pix_240;
		Pix_reg_241 <= Pix_241;
		Pix_reg_242 <= Pix_242;
		Pix_reg_243 <= Pix_243;
		Pix_reg_244 <= Pix_244;
		Pix_reg_245 <= Pix_245;
		Pix_reg_246 <= Pix_246;
		Pix_reg_247 <= Pix_247;
		Pix_reg_248 <= Pix_248;
		Pix_reg_249 <= Pix_249;
		Pix_reg_250 <= Pix_250;
		Pix_reg_251 <= Pix_251;
		Pix_reg_252 <= Pix_252;
		Pix_reg_253 <= Pix_253;
		Pix_reg_254 <= Pix_254;
		Pix_reg_255 <= Pix_255;
		Pix_reg_256 <= Pix_256;
		Pix_reg_257 <= Pix_257;
		Pix_reg_258 <= Pix_258;
		Pix_reg_259 <= Pix_259;
		Pix_reg_260 <= Pix_260;
		Pix_reg_261 <= Pix_261;
		Pix_reg_262 <= Pix_262;
		Pix_reg_263 <= Pix_263;
		Pix_reg_264 <= Pix_264;
		Pix_reg_265 <= Pix_265;
		Pix_reg_266 <= Pix_266;
		Pix_reg_267 <= Pix_267;
		Pix_reg_268 <= Pix_268;
		Pix_reg_269 <= Pix_269;
		Pix_reg_270 <= Pix_270;
		Pix_reg_271 <= Pix_271;
		Pix_reg_272 <= Pix_272;
		Pix_reg_273 <= Pix_273;
		Pix_reg_274 <= Pix_274;
		Pix_reg_275 <= Pix_275;
		Pix_reg_276 <= Pix_276;
		Pix_reg_277 <= Pix_277;
		Pix_reg_278 <= Pix_278;
		Pix_reg_279 <= Pix_279;
		Pix_reg_280 <= Pix_280;
		Pix_reg_281 <= Pix_281;
		Pix_reg_282 <= Pix_282;
		Pix_reg_283 <= Pix_283;
		Pix_reg_284 <= Pix_284;
		Pix_reg_285 <= Pix_285;
		Pix_reg_286 <= Pix_286;
		Pix_reg_287 <= Pix_287;
		Pix_reg_288 <= Pix_288;
		Pix_reg_289 <= Pix_289;
		Pix_reg_290 <= Pix_290;
		Pix_reg_291 <= Pix_291;
		Pix_reg_292 <= Pix_292;
		Pix_reg_293 <= Pix_293;
		Pix_reg_294 <= Pix_294;
		Pix_reg_295 <= Pix_295;
		Pix_reg_296 <= Pix_296;
		Pix_reg_297 <= Pix_297;
		Pix_reg_298 <= Pix_298;
		Pix_reg_299 <= Pix_299;
		Pix_reg_300 <= Pix_300;
		Pix_reg_301 <= Pix_301;
		Pix_reg_302 <= Pix_302;
		Pix_reg_303 <= Pix_303;
		Pix_reg_304 <= Pix_304;
		Pix_reg_305 <= Pix_305;
		Pix_reg_306 <= Pix_306;
		Pix_reg_307 <= Pix_307;
		Pix_reg_308 <= Pix_308;
		Pix_reg_309 <= Pix_309;
		Pix_reg_310 <= Pix_310;
		Pix_reg_311 <= Pix_311;
		Pix_reg_312 <= Pix_312;
		Pix_reg_313 <= Pix_313;
		Pix_reg_314 <= Pix_314;
		Pix_reg_315 <= Pix_315;
		Pix_reg_316 <= Pix_316;
		Pix_reg_317 <= Pix_317;
		Pix_reg_318 <= Pix_318;
		Pix_reg_319 <= Pix_319;
		Pix_reg_320 <= Pix_320;
		Pix_reg_321 <= Pix_321;
		Pix_reg_322 <= Pix_322;
		Pix_reg_323 <= Pix_323;
		Pix_reg_324 <= Pix_324;
		Pix_reg_325 <= Pix_325;
		Pix_reg_326 <= Pix_326;
		Pix_reg_327 <= Pix_327;
		Pix_reg_328 <= Pix_328;
		Pix_reg_329 <= Pix_329;
		Pix_reg_330 <= Pix_330;
		Pix_reg_331 <= Pix_331;
		Pix_reg_332 <= Pix_332;
		Pix_reg_333 <= Pix_333;
		Pix_reg_334 <= Pix_334;
		Pix_reg_335 <= Pix_335;
		Pix_reg_336 <= Pix_336;
		Pix_reg_337 <= Pix_337;
		Pix_reg_338 <= Pix_338;
		Pix_reg_339 <= Pix_339;
		Pix_reg_340 <= Pix_340;
		Pix_reg_341 <= Pix_341;
		Pix_reg_342 <= Pix_342;
		Pix_reg_343 <= Pix_343;
		Pix_reg_344 <= Pix_344;
		Pix_reg_345 <= Pix_345;
		Pix_reg_346 <= Pix_346;
		Pix_reg_347 <= Pix_347;
		Pix_reg_348 <= Pix_348;
		Pix_reg_349 <= Pix_349;
		Pix_reg_350 <= Pix_350;
		Pix_reg_351 <= Pix_351;
		Pix_reg_352 <= Pix_352;
		Pix_reg_353 <= Pix_353;
		Pix_reg_354 <= Pix_354;
		Pix_reg_355 <= Pix_355;
		Pix_reg_356 <= Pix_356;
		Pix_reg_357 <= Pix_357;
		Pix_reg_358 <= Pix_358;
		Pix_reg_359 <= Pix_359;
		Pix_reg_360 <= Pix_360;
		Pix_reg_361 <= Pix_361;
		Pix_reg_362 <= Pix_362;
		Pix_reg_363 <= Pix_363;
		Pix_reg_364 <= Pix_364;
		Pix_reg_365 <= Pix_365;
		Pix_reg_366 <= Pix_366;
		Pix_reg_367 <= Pix_367;
		Pix_reg_368 <= Pix_368;
		Pix_reg_369 <= Pix_369;
		Pix_reg_370 <= Pix_370;
		Pix_reg_371 <= Pix_371;
		Pix_reg_372 <= Pix_372;
		Pix_reg_373 <= Pix_373;
		Pix_reg_374 <= Pix_374;
		Pix_reg_375 <= Pix_375;
		Pix_reg_376 <= Pix_376;
		Pix_reg_377 <= Pix_377;
		Pix_reg_378 <= Pix_378;
		Pix_reg_379 <= Pix_379;
		Pix_reg_380 <= Pix_380;
		Pix_reg_381 <= Pix_381;
		Pix_reg_382 <= Pix_382;
		Pix_reg_383 <= Pix_383;
		Pix_reg_384 <= Pix_384;
		Pix_reg_385 <= Pix_385;
		Pix_reg_386 <= Pix_386;
		Pix_reg_387 <= Pix_387;
		Pix_reg_388 <= Pix_388;
		Pix_reg_389 <= Pix_389;
		Pix_reg_390 <= Pix_390;
		Pix_reg_391 <= Pix_391;
		Pix_reg_392 <= Pix_392;
		Pix_reg_393 <= Pix_393;
		Pix_reg_394 <= Pix_394;
		Pix_reg_395 <= Pix_395;
		Pix_reg_396 <= Pix_396;
		Pix_reg_397 <= Pix_397;
		Pix_reg_398 <= Pix_398;
		Pix_reg_399 <= Pix_399;
		Pix_reg_400 <= Pix_400;
		Pix_reg_401 <= Pix_401;
		Pix_reg_402 <= Pix_402;
		Pix_reg_403 <= Pix_403;
		Pix_reg_404 <= Pix_404;
		Pix_reg_405 <= Pix_405;
		Pix_reg_406 <= Pix_406;
		Pix_reg_407 <= Pix_407;
		Pix_reg_408 <= Pix_408;
		Pix_reg_409 <= Pix_409;
		Pix_reg_410 <= Pix_410;
		Pix_reg_411 <= Pix_411;
		Pix_reg_412 <= Pix_412;
		Pix_reg_413 <= Pix_413;
		Pix_reg_414 <= Pix_414;
		Pix_reg_415 <= Pix_415;
		Pix_reg_416 <= Pix_416;
		Pix_reg_417 <= Pix_417;
		Pix_reg_418 <= Pix_418;
		Pix_reg_419 <= Pix_419;
		Pix_reg_420 <= Pix_420;
		Pix_reg_421 <= Pix_421;
		Pix_reg_422 <= Pix_422;
		Pix_reg_423 <= Pix_423;
		Pix_reg_424 <= Pix_424;
		Pix_reg_425 <= Pix_425;
		Pix_reg_426 <= Pix_426;
		Pix_reg_427 <= Pix_427;
		Pix_reg_428 <= Pix_428;
		Pix_reg_429 <= Pix_429;
		Pix_reg_430 <= Pix_430;
		Pix_reg_431 <= Pix_431;
		Pix_reg_432 <= Pix_432;
		Pix_reg_433 <= Pix_433;
		Pix_reg_434 <= Pix_434;
		Pix_reg_435 <= Pix_435;
		Pix_reg_436 <= Pix_436;
		Pix_reg_437 <= Pix_437;
		Pix_reg_438 <= Pix_438;
		Pix_reg_439 <= Pix_439;
		Pix_reg_440 <= Pix_440;
		Pix_reg_441 <= Pix_441;
		Pix_reg_442 <= Pix_442;
		Pix_reg_443 <= Pix_443;
		Pix_reg_444 <= Pix_444;
		Pix_reg_445 <= Pix_445;
		Pix_reg_446 <= Pix_446;
		Pix_reg_447 <= Pix_447;
		Pix_reg_448 <= Pix_448;
		Pix_reg_449 <= Pix_449;
		Pix_reg_450 <= Pix_450;
		Pix_reg_451 <= Pix_451;
		Pix_reg_452 <= Pix_452;
		Pix_reg_453 <= Pix_453;
		Pix_reg_454 <= Pix_454;
		Pix_reg_455 <= Pix_455;
		Pix_reg_456 <= Pix_456;
		Pix_reg_457 <= Pix_457;
		Pix_reg_458 <= Pix_458;
		Pix_reg_459 <= Pix_459;
		Pix_reg_460 <= Pix_460;
		Pix_reg_461 <= Pix_461;
		Pix_reg_462 <= Pix_462;
		Pix_reg_463 <= Pix_463;
		Pix_reg_464 <= Pix_464;
		Pix_reg_465 <= Pix_465;
		Pix_reg_466 <= Pix_466;
		Pix_reg_467 <= Pix_467;
		Pix_reg_468 <= Pix_468;
		Pix_reg_469 <= Pix_469;
		Pix_reg_470 <= Pix_470;
		Pix_reg_471 <= Pix_471;
		Pix_reg_472 <= Pix_472;
		Pix_reg_473 <= Pix_473;
		Pix_reg_474 <= Pix_474;
		Pix_reg_475 <= Pix_475;
		Pix_reg_476 <= Pix_476;
		Pix_reg_477 <= Pix_477;
		Pix_reg_478 <= Pix_478;
		Pix_reg_479 <= Pix_479;
		Pix_reg_480 <= Pix_480;
		Pix_reg_481 <= Pix_481;
		Pix_reg_482 <= Pix_482;
		Pix_reg_483 <= Pix_483;
		Pix_reg_484 <= Pix_484;
		Pix_reg_485 <= Pix_485;
		Pix_reg_486 <= Pix_486;
		Pix_reg_487 <= Pix_487;
		Pix_reg_488 <= Pix_488;
		Pix_reg_489 <= Pix_489;
		Pix_reg_490 <= Pix_490;
		Pix_reg_491 <= Pix_491;
		Pix_reg_492 <= Pix_492;
		Pix_reg_493 <= Pix_493;
		Pix_reg_494 <= Pix_494;
		Pix_reg_495 <= Pix_495;
		Pix_reg_496 <= Pix_496;
		Pix_reg_497 <= Pix_497;
		Pix_reg_498 <= Pix_498;
		Pix_reg_499 <= Pix_499;
		Pix_reg_500 <= Pix_500;
		Pix_reg_501 <= Pix_501;
		Pix_reg_502 <= Pix_502;
		Pix_reg_503 <= Pix_503;
		Pix_reg_504 <= Pix_504;
		Pix_reg_505 <= Pix_505;
		Pix_reg_506 <= Pix_506;
		Pix_reg_507 <= Pix_507;
		Pix_reg_508 <= Pix_508;
		Pix_reg_509 <= Pix_509;
		Pix_reg_510 <= Pix_510;
		Pix_reg_511 <= Pix_511;
		Pix_reg_512 <= Pix_512;
		Pix_reg_513 <= Pix_513;
		Pix_reg_514 <= Pix_514;
		Pix_reg_515 <= Pix_515;
		Pix_reg_516 <= Pix_516;
		Pix_reg_517 <= Pix_517;
		Pix_reg_518 <= Pix_518;
		Pix_reg_519 <= Pix_519;
		Pix_reg_520 <= Pix_520;
		Pix_reg_521 <= Pix_521;
		Pix_reg_522 <= Pix_522;
		Pix_reg_523 <= Pix_523;
		Pix_reg_524 <= Pix_524;
		Pix_reg_525 <= Pix_525;
		Pix_reg_526 <= Pix_526;
		Pix_reg_527 <= Pix_527;
		Pix_reg_528 <= Pix_528;
		Pix_reg_529 <= Pix_529;
		Pix_reg_530 <= Pix_530;
		Pix_reg_531 <= Pix_531;
		Pix_reg_532 <= Pix_532;
		Pix_reg_533 <= Pix_533;
		Pix_reg_534 <= Pix_534;
		Pix_reg_535 <= Pix_535;
		Pix_reg_536 <= Pix_536;
		Pix_reg_537 <= Pix_537;
		Pix_reg_538 <= Pix_538;
		Pix_reg_539 <= Pix_539;
		Pix_reg_540 <= Pix_540;
		Pix_reg_541 <= Pix_541;
		Pix_reg_542 <= Pix_542;
		Pix_reg_543 <= Pix_543;
		Pix_reg_544 <= Pix_544;
		Pix_reg_545 <= Pix_545;
		Pix_reg_546 <= Pix_546;
		Pix_reg_547 <= Pix_547;
		Pix_reg_548 <= Pix_548;
		Pix_reg_549 <= Pix_549;
		Pix_reg_550 <= Pix_550;
		Pix_reg_551 <= Pix_551;
		Pix_reg_552 <= Pix_552;
		Pix_reg_553 <= Pix_553;
		Pix_reg_554 <= Pix_554;
		Pix_reg_555 <= Pix_555;
		Pix_reg_556 <= Pix_556;
		Pix_reg_557 <= Pix_557;
		Pix_reg_558 <= Pix_558;
		Pix_reg_559 <= Pix_559;
		Pix_reg_560 <= Pix_560;
		Pix_reg_561 <= Pix_561;
		Pix_reg_562 <= Pix_562;
		Pix_reg_563 <= Pix_563;
		Pix_reg_564 <= Pix_564;
		Pix_reg_565 <= Pix_565;
		Pix_reg_566 <= Pix_566;
		Pix_reg_567 <= Pix_567;
		Pix_reg_568 <= Pix_568;
		Pix_reg_569 <= Pix_569;
		Pix_reg_570 <= Pix_570;
		Pix_reg_571 <= Pix_571;
		Pix_reg_572 <= Pix_572;
		Pix_reg_573 <= Pix_573;
		Pix_reg_574 <= Pix_574;
		Pix_reg_575 <= Pix_575;
		Pix_reg_576 <= Pix_576;
		Pix_reg_577 <= Pix_577;
		Pix_reg_578 <= Pix_578;
		Pix_reg_579 <= Pix_579;
		Pix_reg_580 <= Pix_580;
		Pix_reg_581 <= Pix_581;
		Pix_reg_582 <= Pix_582;
		Pix_reg_583 <= Pix_583;
		Pix_reg_584 <= Pix_584;
		Pix_reg_585 <= Pix_585;
		Pix_reg_586 <= Pix_586;
		Pix_reg_587 <= Pix_587;
		Pix_reg_588 <= Pix_588;
		Pix_reg_589 <= Pix_589;
		Pix_reg_590 <= Pix_590;
		Pix_reg_591 <= Pix_591;
		Pix_reg_592 <= Pix_592;
		Pix_reg_593 <= Pix_593;
		Pix_reg_594 <= Pix_594;
		Pix_reg_595 <= Pix_595;
		Pix_reg_596 <= Pix_596;
		Pix_reg_597 <= Pix_597;
		Pix_reg_598 <= Pix_598;
		Pix_reg_599 <= Pix_599;
		Pix_reg_600 <= Pix_600;
		Pix_reg_601 <= Pix_601;
		Pix_reg_602 <= Pix_602;
		Pix_reg_603 <= Pix_603;
		Pix_reg_604 <= Pix_604;
		Pix_reg_605 <= Pix_605;
		Pix_reg_606 <= Pix_606;
		Pix_reg_607 <= Pix_607;
		Pix_reg_608 <= Pix_608;
		Pix_reg_609 <= Pix_609;
		Pix_reg_610 <= Pix_610;
		Pix_reg_611 <= Pix_611;
		Pix_reg_612 <= Pix_612;
		Pix_reg_613 <= Pix_613;
		Pix_reg_614 <= Pix_614;
		Pix_reg_615 <= Pix_615;
		Pix_reg_616 <= Pix_616;
		Pix_reg_617 <= Pix_617;
		Pix_reg_618 <= Pix_618;
		Pix_reg_619 <= Pix_619;
		Pix_reg_620 <= Pix_620;
		Pix_reg_621 <= Pix_621;
		Pix_reg_622 <= Pix_622;
		Pix_reg_623 <= Pix_623;
		Pix_reg_624 <= Pix_624;
		Pix_reg_625 <= Pix_625;
		Pix_reg_626 <= Pix_626;
		Pix_reg_627 <= Pix_627;
		Pix_reg_628 <= Pix_628;
		Pix_reg_629 <= Pix_629;
		Pix_reg_630 <= Pix_630;
		Pix_reg_631 <= Pix_631;
		Pix_reg_632 <= Pix_632;
		Pix_reg_633 <= Pix_633;
		Pix_reg_634 <= Pix_634;
		Pix_reg_635 <= Pix_635;
		Pix_reg_636 <= Pix_636;
		Pix_reg_637 <= Pix_637;
		Pix_reg_638 <= Pix_638;
		Pix_reg_639 <= Pix_639;
		Pix_reg_640 <= Pix_640;
		Pix_reg_641 <= Pix_641;
		Pix_reg_642 <= Pix_642;
		Pix_reg_643 <= Pix_643;
		Pix_reg_644 <= Pix_644;
		Pix_reg_645 <= Pix_645;
		Pix_reg_646 <= Pix_646;
		Pix_reg_647 <= Pix_647;
		Pix_reg_648 <= Pix_648;
		Pix_reg_649 <= Pix_649;
		Pix_reg_650 <= Pix_650;
		Pix_reg_651 <= Pix_651;
		Pix_reg_652 <= Pix_652;
		Pix_reg_653 <= Pix_653;
		Pix_reg_654 <= Pix_654;
		Pix_reg_655 <= Pix_655;
		Pix_reg_656 <= Pix_656;
		Pix_reg_657 <= Pix_657;
		Pix_reg_658 <= Pix_658;
		Pix_reg_659 <= Pix_659;
		Pix_reg_660 <= Pix_660;
		Pix_reg_661 <= Pix_661;
		Pix_reg_662 <= Pix_662;
		Pix_reg_663 <= Pix_663;
		Pix_reg_664 <= Pix_664;
		Pix_reg_665 <= Pix_665;
		Pix_reg_666 <= Pix_666;
		Pix_reg_667 <= Pix_667;
		Pix_reg_668 <= Pix_668;
		Pix_reg_669 <= Pix_669;
		Pix_reg_670 <= Pix_670;
		Pix_reg_671 <= Pix_671;
		Pix_reg_672 <= Pix_672;
		Pix_reg_673 <= Pix_673;
		Pix_reg_674 <= Pix_674;
		Pix_reg_675 <= Pix_675;
		Pix_reg_676 <= Pix_676;
		Pix_reg_677 <= Pix_677;
		Pix_reg_678 <= Pix_678;
		Pix_reg_679 <= Pix_679;
		Pix_reg_680 <= Pix_680;
		Pix_reg_681 <= Pix_681;
		Pix_reg_682 <= Pix_682;
		Pix_reg_683 <= Pix_683;
		Pix_reg_684 <= Pix_684;
		Pix_reg_685 <= Pix_685;
		Pix_reg_686 <= Pix_686;
		Pix_reg_687 <= Pix_687;
		Pix_reg_688 <= Pix_688;
		Pix_reg_689 <= Pix_689;
		Pix_reg_690 <= Pix_690;
		Pix_reg_691 <= Pix_691;
		Pix_reg_692 <= Pix_692;
		Pix_reg_693 <= Pix_693;
		Pix_reg_694 <= Pix_694;
		Pix_reg_695 <= Pix_695;
		Pix_reg_696 <= Pix_696;
		Pix_reg_697 <= Pix_697;
		Pix_reg_698 <= Pix_698;
		Pix_reg_699 <= Pix_699;
		Pix_reg_700 <= Pix_700;
		Pix_reg_701 <= Pix_701;
		Pix_reg_702 <= Pix_702;
		Pix_reg_703 <= Pix_703;
		Pix_reg_704 <= Pix_704;
		Pix_reg_705 <= Pix_705;
		Pix_reg_706 <= Pix_706;
		Pix_reg_707 <= Pix_707;
		Pix_reg_708 <= Pix_708;
		Pix_reg_709 <= Pix_709;
		Pix_reg_710 <= Pix_710;
		Pix_reg_711 <= Pix_711;
		Pix_reg_712 <= Pix_712;
		Pix_reg_713 <= Pix_713;
		Pix_reg_714 <= Pix_714;
		Pix_reg_715 <= Pix_715;
		Pix_reg_716 <= Pix_716;
		Pix_reg_717 <= Pix_717;
		Pix_reg_718 <= Pix_718;
		Pix_reg_719 <= Pix_719;
		Pix_reg_720 <= Pix_720;
		Pix_reg_721 <= Pix_721;
		Pix_reg_722 <= Pix_722;
		Pix_reg_723 <= Pix_723;
		Pix_reg_724 <= Pix_724;
		Pix_reg_725 <= Pix_725;
		Pix_reg_726 <= Pix_726;
		Pix_reg_727 <= Pix_727;
		Pix_reg_728 <= Pix_728;
		Pix_reg_729 <= Pix_729;
		Pix_reg_730 <= Pix_730;
		Pix_reg_731 <= Pix_731;
		Pix_reg_732 <= Pix_732;
		Pix_reg_733 <= Pix_733;
		Pix_reg_734 <= Pix_734;
		Pix_reg_735 <= Pix_735;
		Pix_reg_736 <= Pix_736;
		Pix_reg_737 <= Pix_737;
		Pix_reg_738 <= Pix_738;
		Pix_reg_739 <= Pix_739;
		Pix_reg_740 <= Pix_740;
		Pix_reg_741 <= Pix_741;
		Pix_reg_742 <= Pix_742;
		Pix_reg_743 <= Pix_743;
		Pix_reg_744 <= Pix_744;
		Pix_reg_745 <= Pix_745;
		Pix_reg_746 <= Pix_746;
		Pix_reg_747 <= Pix_747;
		Pix_reg_748 <= Pix_748;
		Pix_reg_749 <= Pix_749;
		Pix_reg_750 <= Pix_750;
		Pix_reg_751 <= Pix_751;
		Pix_reg_752 <= Pix_752;
		Pix_reg_753 <= Pix_753;
		Pix_reg_754 <= Pix_754;
		Pix_reg_755 <= Pix_755;
		Pix_reg_756 <= Pix_756;
		Pix_reg_757 <= Pix_757;
		Pix_reg_758 <= Pix_758;
		Pix_reg_759 <= Pix_759;
		Pix_reg_760 <= Pix_760;
		Pix_reg_761 <= Pix_761;
		Pix_reg_762 <= Pix_762;
		Pix_reg_763 <= Pix_763;
		Pix_reg_764 <= Pix_764;
		Pix_reg_765 <= Pix_765;
		Pix_reg_766 <= Pix_766;
		Pix_reg_767 <= Pix_767;
		Pix_reg_768 <= Pix_768;
		Pix_reg_769 <= Pix_769;
		Pix_reg_770 <= Pix_770;
		Pix_reg_771 <= Pix_771;
		Pix_reg_772 <= Pix_772;
		Pix_reg_773 <= Pix_773;
		Pix_reg_774 <= Pix_774;
		Pix_reg_775 <= Pix_775;
		Pix_reg_776 <= Pix_776;
		Pix_reg_777 <= Pix_777;
		Pix_reg_778 <= Pix_778;
		Pix_reg_779 <= Pix_779;
		Pix_reg_780 <= Pix_780;
		Pix_reg_781 <= Pix_781;
		Pix_reg_782 <= Pix_782;
		Pix_reg_783 <= Pix_783;
		Pix_reg_784 <= Pix_784;

		Wgt_reg_0 <= Wgt_0;
		Wgt_reg_1 <= Wgt_1;
		Wgt_reg_2 <= Wgt_2;
		Wgt_reg_3 <= Wgt_3;
		Wgt_reg_4 <= Wgt_4;
		Wgt_reg_5 <= Wgt_5;
		Wgt_reg_6 <= Wgt_6;
		Wgt_reg_7 <= Wgt_7;
		Wgt_reg_8 <= Wgt_8;
		Wgt_reg_9 <= Wgt_9;
		Wgt_reg_10 <= Wgt_10;
		Wgt_reg_11 <= Wgt_11;
		Wgt_reg_12 <= Wgt_12;
		Wgt_reg_13 <= Wgt_13;
		Wgt_reg_14 <= Wgt_14;
		Wgt_reg_15 <= Wgt_15;
		Wgt_reg_16 <= Wgt_16;
		Wgt_reg_17 <= Wgt_17;
		Wgt_reg_18 <= Wgt_18;
		Wgt_reg_19 <= Wgt_19;
		Wgt_reg_20 <= Wgt_20;
		Wgt_reg_21 <= Wgt_21;
		Wgt_reg_22 <= Wgt_22;
		Wgt_reg_23 <= Wgt_23;
		Wgt_reg_24 <= Wgt_24;
		Wgt_reg_25 <= Wgt_25;
		Wgt_reg_26 <= Wgt_26;
		Wgt_reg_27 <= Wgt_27;
		Wgt_reg_28 <= Wgt_28;
		Wgt_reg_29 <= Wgt_29;
		Wgt_reg_30 <= Wgt_30;
		Wgt_reg_31 <= Wgt_31;
		Wgt_reg_32 <= Wgt_32;
		Wgt_reg_33 <= Wgt_33;
		Wgt_reg_34 <= Wgt_34;
		Wgt_reg_35 <= Wgt_35;
		Wgt_reg_36 <= Wgt_36;
		Wgt_reg_37 <= Wgt_37;
		Wgt_reg_38 <= Wgt_38;
		Wgt_reg_39 <= Wgt_39;
		Wgt_reg_40 <= Wgt_40;
		Wgt_reg_41 <= Wgt_41;
		Wgt_reg_42 <= Wgt_42;
		Wgt_reg_43 <= Wgt_43;
		Wgt_reg_44 <= Wgt_44;
		Wgt_reg_45 <= Wgt_45;
		Wgt_reg_46 <= Wgt_46;
		Wgt_reg_47 <= Wgt_47;
		Wgt_reg_48 <= Wgt_48;
		Wgt_reg_49 <= Wgt_49;
		Wgt_reg_50 <= Wgt_50;
		Wgt_reg_51 <= Wgt_51;
		Wgt_reg_52 <= Wgt_52;
		Wgt_reg_53 <= Wgt_53;
		Wgt_reg_54 <= Wgt_54;
		Wgt_reg_55 <= Wgt_55;
		Wgt_reg_56 <= Wgt_56;
		Wgt_reg_57 <= Wgt_57;
		Wgt_reg_58 <= Wgt_58;
		Wgt_reg_59 <= Wgt_59;
		Wgt_reg_60 <= Wgt_60;
		Wgt_reg_61 <= Wgt_61;
		Wgt_reg_62 <= Wgt_62;
		Wgt_reg_63 <= Wgt_63;
		Wgt_reg_64 <= Wgt_64;
		Wgt_reg_65 <= Wgt_65;
		Wgt_reg_66 <= Wgt_66;
		Wgt_reg_67 <= Wgt_67;
		Wgt_reg_68 <= Wgt_68;
		Wgt_reg_69 <= Wgt_69;
		Wgt_reg_70 <= Wgt_70;
		Wgt_reg_71 <= Wgt_71;
		Wgt_reg_72 <= Wgt_72;
		Wgt_reg_73 <= Wgt_73;
		Wgt_reg_74 <= Wgt_74;
		Wgt_reg_75 <= Wgt_75;
		Wgt_reg_76 <= Wgt_76;
		Wgt_reg_77 <= Wgt_77;
		Wgt_reg_78 <= Wgt_78;
		Wgt_reg_79 <= Wgt_79;
		Wgt_reg_80 <= Wgt_80;
		Wgt_reg_81 <= Wgt_81;
		Wgt_reg_82 <= Wgt_82;
		Wgt_reg_83 <= Wgt_83;
		Wgt_reg_84 <= Wgt_84;
		Wgt_reg_85 <= Wgt_85;
		Wgt_reg_86 <= Wgt_86;
		Wgt_reg_87 <= Wgt_87;
		Wgt_reg_88 <= Wgt_88;
		Wgt_reg_89 <= Wgt_89;
		Wgt_reg_90 <= Wgt_90;
		Wgt_reg_91 <= Wgt_91;
		Wgt_reg_92 <= Wgt_92;
		Wgt_reg_93 <= Wgt_93;
		Wgt_reg_94 <= Wgt_94;
		Wgt_reg_95 <= Wgt_95;
		Wgt_reg_96 <= Wgt_96;
		Wgt_reg_97 <= Wgt_97;
		Wgt_reg_98 <= Wgt_98;
		Wgt_reg_99 <= Wgt_99;
		Wgt_reg_100 <= Wgt_100;
		Wgt_reg_101 <= Wgt_101;
		Wgt_reg_102 <= Wgt_102;
		Wgt_reg_103 <= Wgt_103;
		Wgt_reg_104 <= Wgt_104;
		Wgt_reg_105 <= Wgt_105;
		Wgt_reg_106 <= Wgt_106;
		Wgt_reg_107 <= Wgt_107;
		Wgt_reg_108 <= Wgt_108;
		Wgt_reg_109 <= Wgt_109;
		Wgt_reg_110 <= Wgt_110;
		Wgt_reg_111 <= Wgt_111;
		Wgt_reg_112 <= Wgt_112;
		Wgt_reg_113 <= Wgt_113;
		Wgt_reg_114 <= Wgt_114;
		Wgt_reg_115 <= Wgt_115;
		Wgt_reg_116 <= Wgt_116;
		Wgt_reg_117 <= Wgt_117;
		Wgt_reg_118 <= Wgt_118;
		Wgt_reg_119 <= Wgt_119;
		Wgt_reg_120 <= Wgt_120;
		Wgt_reg_121 <= Wgt_121;
		Wgt_reg_122 <= Wgt_122;
		Wgt_reg_123 <= Wgt_123;
		Wgt_reg_124 <= Wgt_124;
		Wgt_reg_125 <= Wgt_125;
		Wgt_reg_126 <= Wgt_126;
		Wgt_reg_127 <= Wgt_127;
		Wgt_reg_128 <= Wgt_128;
		Wgt_reg_129 <= Wgt_129;
		Wgt_reg_130 <= Wgt_130;
		Wgt_reg_131 <= Wgt_131;
		Wgt_reg_132 <= Wgt_132;
		Wgt_reg_133 <= Wgt_133;
		Wgt_reg_134 <= Wgt_134;
		Wgt_reg_135 <= Wgt_135;
		Wgt_reg_136 <= Wgt_136;
		Wgt_reg_137 <= Wgt_137;
		Wgt_reg_138 <= Wgt_138;
		Wgt_reg_139 <= Wgt_139;
		Wgt_reg_140 <= Wgt_140;
		Wgt_reg_141 <= Wgt_141;
		Wgt_reg_142 <= Wgt_142;
		Wgt_reg_143 <= Wgt_143;
		Wgt_reg_144 <= Wgt_144;
		Wgt_reg_145 <= Wgt_145;
		Wgt_reg_146 <= Wgt_146;
		Wgt_reg_147 <= Wgt_147;
		Wgt_reg_148 <= Wgt_148;
		Wgt_reg_149 <= Wgt_149;
		Wgt_reg_150 <= Wgt_150;
		Wgt_reg_151 <= Wgt_151;
		Wgt_reg_152 <= Wgt_152;
		Wgt_reg_153 <= Wgt_153;
		Wgt_reg_154 <= Wgt_154;
		Wgt_reg_155 <= Wgt_155;
		Wgt_reg_156 <= Wgt_156;
		Wgt_reg_157 <= Wgt_157;
		Wgt_reg_158 <= Wgt_158;
		Wgt_reg_159 <= Wgt_159;
		Wgt_reg_160 <= Wgt_160;
		Wgt_reg_161 <= Wgt_161;
		Wgt_reg_162 <= Wgt_162;
		Wgt_reg_163 <= Wgt_163;
		Wgt_reg_164 <= Wgt_164;
		Wgt_reg_165 <= Wgt_165;
		Wgt_reg_166 <= Wgt_166;
		Wgt_reg_167 <= Wgt_167;
		Wgt_reg_168 <= Wgt_168;
		Wgt_reg_169 <= Wgt_169;
		Wgt_reg_170 <= Wgt_170;
		Wgt_reg_171 <= Wgt_171;
		Wgt_reg_172 <= Wgt_172;
		Wgt_reg_173 <= Wgt_173;
		Wgt_reg_174 <= Wgt_174;
		Wgt_reg_175 <= Wgt_175;
		Wgt_reg_176 <= Wgt_176;
		Wgt_reg_177 <= Wgt_177;
		Wgt_reg_178 <= Wgt_178;
		Wgt_reg_179 <= Wgt_179;
		Wgt_reg_180 <= Wgt_180;
		Wgt_reg_181 <= Wgt_181;
		Wgt_reg_182 <= Wgt_182;
		Wgt_reg_183 <= Wgt_183;
		Wgt_reg_184 <= Wgt_184;
		Wgt_reg_185 <= Wgt_185;
		Wgt_reg_186 <= Wgt_186;
		Wgt_reg_187 <= Wgt_187;
		Wgt_reg_188 <= Wgt_188;
		Wgt_reg_189 <= Wgt_189;
		Wgt_reg_190 <= Wgt_190;
		Wgt_reg_191 <= Wgt_191;
		Wgt_reg_192 <= Wgt_192;
		Wgt_reg_193 <= Wgt_193;
		Wgt_reg_194 <= Wgt_194;
		Wgt_reg_195 <= Wgt_195;
		Wgt_reg_196 <= Wgt_196;
		Wgt_reg_197 <= Wgt_197;
		Wgt_reg_198 <= Wgt_198;
		Wgt_reg_199 <= Wgt_199;
		Wgt_reg_200 <= Wgt_200;
		Wgt_reg_201 <= Wgt_201;
		Wgt_reg_202 <= Wgt_202;
		Wgt_reg_203 <= Wgt_203;
		Wgt_reg_204 <= Wgt_204;
		Wgt_reg_205 <= Wgt_205;
		Wgt_reg_206 <= Wgt_206;
		Wgt_reg_207 <= Wgt_207;
		Wgt_reg_208 <= Wgt_208;
		Wgt_reg_209 <= Wgt_209;
		Wgt_reg_210 <= Wgt_210;
		Wgt_reg_211 <= Wgt_211;
		Wgt_reg_212 <= Wgt_212;
		Wgt_reg_213 <= Wgt_213;
		Wgt_reg_214 <= Wgt_214;
		Wgt_reg_215 <= Wgt_215;
		Wgt_reg_216 <= Wgt_216;
		Wgt_reg_217 <= Wgt_217;
		Wgt_reg_218 <= Wgt_218;
		Wgt_reg_219 <= Wgt_219;
		Wgt_reg_220 <= Wgt_220;
		Wgt_reg_221 <= Wgt_221;
		Wgt_reg_222 <= Wgt_222;
		Wgt_reg_223 <= Wgt_223;
		Wgt_reg_224 <= Wgt_224;
		Wgt_reg_225 <= Wgt_225;
		Wgt_reg_226 <= Wgt_226;
		Wgt_reg_227 <= Wgt_227;
		Wgt_reg_228 <= Wgt_228;
		Wgt_reg_229 <= Wgt_229;
		Wgt_reg_230 <= Wgt_230;
		Wgt_reg_231 <= Wgt_231;
		Wgt_reg_232 <= Wgt_232;
		Wgt_reg_233 <= Wgt_233;
		Wgt_reg_234 <= Wgt_234;
		Wgt_reg_235 <= Wgt_235;
		Wgt_reg_236 <= Wgt_236;
		Wgt_reg_237 <= Wgt_237;
		Wgt_reg_238 <= Wgt_238;
		Wgt_reg_239 <= Wgt_239;
		Wgt_reg_240 <= Wgt_240;
		Wgt_reg_241 <= Wgt_241;
		Wgt_reg_242 <= Wgt_242;
		Wgt_reg_243 <= Wgt_243;
		Wgt_reg_244 <= Wgt_244;
		Wgt_reg_245 <= Wgt_245;
		Wgt_reg_246 <= Wgt_246;
		Wgt_reg_247 <= Wgt_247;
		Wgt_reg_248 <= Wgt_248;
		Wgt_reg_249 <= Wgt_249;
		Wgt_reg_250 <= Wgt_250;
		Wgt_reg_251 <= Wgt_251;
		Wgt_reg_252 <= Wgt_252;
		Wgt_reg_253 <= Wgt_253;
		Wgt_reg_254 <= Wgt_254;
		Wgt_reg_255 <= Wgt_255;
		Wgt_reg_256 <= Wgt_256;
		Wgt_reg_257 <= Wgt_257;
		Wgt_reg_258 <= Wgt_258;
		Wgt_reg_259 <= Wgt_259;
		Wgt_reg_260 <= Wgt_260;
		Wgt_reg_261 <= Wgt_261;
		Wgt_reg_262 <= Wgt_262;
		Wgt_reg_263 <= Wgt_263;
		Wgt_reg_264 <= Wgt_264;
		Wgt_reg_265 <= Wgt_265;
		Wgt_reg_266 <= Wgt_266;
		Wgt_reg_267 <= Wgt_267;
		Wgt_reg_268 <= Wgt_268;
		Wgt_reg_269 <= Wgt_269;
		Wgt_reg_270 <= Wgt_270;
		Wgt_reg_271 <= Wgt_271;
		Wgt_reg_272 <= Wgt_272;
		Wgt_reg_273 <= Wgt_273;
		Wgt_reg_274 <= Wgt_274;
		Wgt_reg_275 <= Wgt_275;
		Wgt_reg_276 <= Wgt_276;
		Wgt_reg_277 <= Wgt_277;
		Wgt_reg_278 <= Wgt_278;
		Wgt_reg_279 <= Wgt_279;
		Wgt_reg_280 <= Wgt_280;
		Wgt_reg_281 <= Wgt_281;
		Wgt_reg_282 <= Wgt_282;
		Wgt_reg_283 <= Wgt_283;
		Wgt_reg_284 <= Wgt_284;
		Wgt_reg_285 <= Wgt_285;
		Wgt_reg_286 <= Wgt_286;
		Wgt_reg_287 <= Wgt_287;
		Wgt_reg_288 <= Wgt_288;
		Wgt_reg_289 <= Wgt_289;
		Wgt_reg_290 <= Wgt_290;
		Wgt_reg_291 <= Wgt_291;
		Wgt_reg_292 <= Wgt_292;
		Wgt_reg_293 <= Wgt_293;
		Wgt_reg_294 <= Wgt_294;
		Wgt_reg_295 <= Wgt_295;
		Wgt_reg_296 <= Wgt_296;
		Wgt_reg_297 <= Wgt_297;
		Wgt_reg_298 <= Wgt_298;
		Wgt_reg_299 <= Wgt_299;
		Wgt_reg_300 <= Wgt_300;
		Wgt_reg_301 <= Wgt_301;
		Wgt_reg_302 <= Wgt_302;
		Wgt_reg_303 <= Wgt_303;
		Wgt_reg_304 <= Wgt_304;
		Wgt_reg_305 <= Wgt_305;
		Wgt_reg_306 <= Wgt_306;
		Wgt_reg_307 <= Wgt_307;
		Wgt_reg_308 <= Wgt_308;
		Wgt_reg_309 <= Wgt_309;
		Wgt_reg_310 <= Wgt_310;
		Wgt_reg_311 <= Wgt_311;
		Wgt_reg_312 <= Wgt_312;
		Wgt_reg_313 <= Wgt_313;
		Wgt_reg_314 <= Wgt_314;
		Wgt_reg_315 <= Wgt_315;
		Wgt_reg_316 <= Wgt_316;
		Wgt_reg_317 <= Wgt_317;
		Wgt_reg_318 <= Wgt_318;
		Wgt_reg_319 <= Wgt_319;
		Wgt_reg_320 <= Wgt_320;
		Wgt_reg_321 <= Wgt_321;
		Wgt_reg_322 <= Wgt_322;
		Wgt_reg_323 <= Wgt_323;
		Wgt_reg_324 <= Wgt_324;
		Wgt_reg_325 <= Wgt_325;
		Wgt_reg_326 <= Wgt_326;
		Wgt_reg_327 <= Wgt_327;
		Wgt_reg_328 <= Wgt_328;
		Wgt_reg_329 <= Wgt_329;
		Wgt_reg_330 <= Wgt_330;
		Wgt_reg_331 <= Wgt_331;
		Wgt_reg_332 <= Wgt_332;
		Wgt_reg_333 <= Wgt_333;
		Wgt_reg_334 <= Wgt_334;
		Wgt_reg_335 <= Wgt_335;
		Wgt_reg_336 <= Wgt_336;
		Wgt_reg_337 <= Wgt_337;
		Wgt_reg_338 <= Wgt_338;
		Wgt_reg_339 <= Wgt_339;
		Wgt_reg_340 <= Wgt_340;
		Wgt_reg_341 <= Wgt_341;
		Wgt_reg_342 <= Wgt_342;
		Wgt_reg_343 <= Wgt_343;
		Wgt_reg_344 <= Wgt_344;
		Wgt_reg_345 <= Wgt_345;
		Wgt_reg_346 <= Wgt_346;
		Wgt_reg_347 <= Wgt_347;
		Wgt_reg_348 <= Wgt_348;
		Wgt_reg_349 <= Wgt_349;
		Wgt_reg_350 <= Wgt_350;
		Wgt_reg_351 <= Wgt_351;
		Wgt_reg_352 <= Wgt_352;
		Wgt_reg_353 <= Wgt_353;
		Wgt_reg_354 <= Wgt_354;
		Wgt_reg_355 <= Wgt_355;
		Wgt_reg_356 <= Wgt_356;
		Wgt_reg_357 <= Wgt_357;
		Wgt_reg_358 <= Wgt_358;
		Wgt_reg_359 <= Wgt_359;
		Wgt_reg_360 <= Wgt_360;
		Wgt_reg_361 <= Wgt_361;
		Wgt_reg_362 <= Wgt_362;
		Wgt_reg_363 <= Wgt_363;
		Wgt_reg_364 <= Wgt_364;
		Wgt_reg_365 <= Wgt_365;
		Wgt_reg_366 <= Wgt_366;
		Wgt_reg_367 <= Wgt_367;
		Wgt_reg_368 <= Wgt_368;
		Wgt_reg_369 <= Wgt_369;
		Wgt_reg_370 <= Wgt_370;
		Wgt_reg_371 <= Wgt_371;
		Wgt_reg_372 <= Wgt_372;
		Wgt_reg_373 <= Wgt_373;
		Wgt_reg_374 <= Wgt_374;
		Wgt_reg_375 <= Wgt_375;
		Wgt_reg_376 <= Wgt_376;
		Wgt_reg_377 <= Wgt_377;
		Wgt_reg_378 <= Wgt_378;
		Wgt_reg_379 <= Wgt_379;
		Wgt_reg_380 <= Wgt_380;
		Wgt_reg_381 <= Wgt_381;
		Wgt_reg_382 <= Wgt_382;
		Wgt_reg_383 <= Wgt_383;
		Wgt_reg_384 <= Wgt_384;
		Wgt_reg_385 <= Wgt_385;
		Wgt_reg_386 <= Wgt_386;
		Wgt_reg_387 <= Wgt_387;
		Wgt_reg_388 <= Wgt_388;
		Wgt_reg_389 <= Wgt_389;
		Wgt_reg_390 <= Wgt_390;
		Wgt_reg_391 <= Wgt_391;
		Wgt_reg_392 <= Wgt_392;
		Wgt_reg_393 <= Wgt_393;
		Wgt_reg_394 <= Wgt_394;
		Wgt_reg_395 <= Wgt_395;
		Wgt_reg_396 <= Wgt_396;
		Wgt_reg_397 <= Wgt_397;
		Wgt_reg_398 <= Wgt_398;
		Wgt_reg_399 <= Wgt_399;
		Wgt_reg_400 <= Wgt_400;
		Wgt_reg_401 <= Wgt_401;
		Wgt_reg_402 <= Wgt_402;
		Wgt_reg_403 <= Wgt_403;
		Wgt_reg_404 <= Wgt_404;
		Wgt_reg_405 <= Wgt_405;
		Wgt_reg_406 <= Wgt_406;
		Wgt_reg_407 <= Wgt_407;
		Wgt_reg_408 <= Wgt_408;
		Wgt_reg_409 <= Wgt_409;
		Wgt_reg_410 <= Wgt_410;
		Wgt_reg_411 <= Wgt_411;
		Wgt_reg_412 <= Wgt_412;
		Wgt_reg_413 <= Wgt_413;
		Wgt_reg_414 <= Wgt_414;
		Wgt_reg_415 <= Wgt_415;
		Wgt_reg_416 <= Wgt_416;
		Wgt_reg_417 <= Wgt_417;
		Wgt_reg_418 <= Wgt_418;
		Wgt_reg_419 <= Wgt_419;
		Wgt_reg_420 <= Wgt_420;
		Wgt_reg_421 <= Wgt_421;
		Wgt_reg_422 <= Wgt_422;
		Wgt_reg_423 <= Wgt_423;
		Wgt_reg_424 <= Wgt_424;
		Wgt_reg_425 <= Wgt_425;
		Wgt_reg_426 <= Wgt_426;
		Wgt_reg_427 <= Wgt_427;
		Wgt_reg_428 <= Wgt_428;
		Wgt_reg_429 <= Wgt_429;
		Wgt_reg_430 <= Wgt_430;
		Wgt_reg_431 <= Wgt_431;
		Wgt_reg_432 <= Wgt_432;
		Wgt_reg_433 <= Wgt_433;
		Wgt_reg_434 <= Wgt_434;
		Wgt_reg_435 <= Wgt_435;
		Wgt_reg_436 <= Wgt_436;
		Wgt_reg_437 <= Wgt_437;
		Wgt_reg_438 <= Wgt_438;
		Wgt_reg_439 <= Wgt_439;
		Wgt_reg_440 <= Wgt_440;
		Wgt_reg_441 <= Wgt_441;
		Wgt_reg_442 <= Wgt_442;
		Wgt_reg_443 <= Wgt_443;
		Wgt_reg_444 <= Wgt_444;
		Wgt_reg_445 <= Wgt_445;
		Wgt_reg_446 <= Wgt_446;
		Wgt_reg_447 <= Wgt_447;
		Wgt_reg_448 <= Wgt_448;
		Wgt_reg_449 <= Wgt_449;
		Wgt_reg_450 <= Wgt_450;
		Wgt_reg_451 <= Wgt_451;
		Wgt_reg_452 <= Wgt_452;
		Wgt_reg_453 <= Wgt_453;
		Wgt_reg_454 <= Wgt_454;
		Wgt_reg_455 <= Wgt_455;
		Wgt_reg_456 <= Wgt_456;
		Wgt_reg_457 <= Wgt_457;
		Wgt_reg_458 <= Wgt_458;
		Wgt_reg_459 <= Wgt_459;
		Wgt_reg_460 <= Wgt_460;
		Wgt_reg_461 <= Wgt_461;
		Wgt_reg_462 <= Wgt_462;
		Wgt_reg_463 <= Wgt_463;
		Wgt_reg_464 <= Wgt_464;
		Wgt_reg_465 <= Wgt_465;
		Wgt_reg_466 <= Wgt_466;
		Wgt_reg_467 <= Wgt_467;
		Wgt_reg_468 <= Wgt_468;
		Wgt_reg_469 <= Wgt_469;
		Wgt_reg_470 <= Wgt_470;
		Wgt_reg_471 <= Wgt_471;
		Wgt_reg_472 <= Wgt_472;
		Wgt_reg_473 <= Wgt_473;
		Wgt_reg_474 <= Wgt_474;
		Wgt_reg_475 <= Wgt_475;
		Wgt_reg_476 <= Wgt_476;
		Wgt_reg_477 <= Wgt_477;
		Wgt_reg_478 <= Wgt_478;
		Wgt_reg_479 <= Wgt_479;
		Wgt_reg_480 <= Wgt_480;
		Wgt_reg_481 <= Wgt_481;
		Wgt_reg_482 <= Wgt_482;
		Wgt_reg_483 <= Wgt_483;
		Wgt_reg_484 <= Wgt_484;
		Wgt_reg_485 <= Wgt_485;
		Wgt_reg_486 <= Wgt_486;
		Wgt_reg_487 <= Wgt_487;
		Wgt_reg_488 <= Wgt_488;
		Wgt_reg_489 <= Wgt_489;
		Wgt_reg_490 <= Wgt_490;
		Wgt_reg_491 <= Wgt_491;
		Wgt_reg_492 <= Wgt_492;
		Wgt_reg_493 <= Wgt_493;
		Wgt_reg_494 <= Wgt_494;
		Wgt_reg_495 <= Wgt_495;
		Wgt_reg_496 <= Wgt_496;
		Wgt_reg_497 <= Wgt_497;
		Wgt_reg_498 <= Wgt_498;
		Wgt_reg_499 <= Wgt_499;
		Wgt_reg_500 <= Wgt_500;
		Wgt_reg_501 <= Wgt_501;
		Wgt_reg_502 <= Wgt_502;
		Wgt_reg_503 <= Wgt_503;
		Wgt_reg_504 <= Wgt_504;
		Wgt_reg_505 <= Wgt_505;
		Wgt_reg_506 <= Wgt_506;
		Wgt_reg_507 <= Wgt_507;
		Wgt_reg_508 <= Wgt_508;
		Wgt_reg_509 <= Wgt_509;
		Wgt_reg_510 <= Wgt_510;
		Wgt_reg_511 <= Wgt_511;
		Wgt_reg_512 <= Wgt_512;
		Wgt_reg_513 <= Wgt_513;
		Wgt_reg_514 <= Wgt_514;
		Wgt_reg_515 <= Wgt_515;
		Wgt_reg_516 <= Wgt_516;
		Wgt_reg_517 <= Wgt_517;
		Wgt_reg_518 <= Wgt_518;
		Wgt_reg_519 <= Wgt_519;
		Wgt_reg_520 <= Wgt_520;
		Wgt_reg_521 <= Wgt_521;
		Wgt_reg_522 <= Wgt_522;
		Wgt_reg_523 <= Wgt_523;
		Wgt_reg_524 <= Wgt_524;
		Wgt_reg_525 <= Wgt_525;
		Wgt_reg_526 <= Wgt_526;
		Wgt_reg_527 <= Wgt_527;
		Wgt_reg_528 <= Wgt_528;
		Wgt_reg_529 <= Wgt_529;
		Wgt_reg_530 <= Wgt_530;
		Wgt_reg_531 <= Wgt_531;
		Wgt_reg_532 <= Wgt_532;
		Wgt_reg_533 <= Wgt_533;
		Wgt_reg_534 <= Wgt_534;
		Wgt_reg_535 <= Wgt_535;
		Wgt_reg_536 <= Wgt_536;
		Wgt_reg_537 <= Wgt_537;
		Wgt_reg_538 <= Wgt_538;
		Wgt_reg_539 <= Wgt_539;
		Wgt_reg_540 <= Wgt_540;
		Wgt_reg_541 <= Wgt_541;
		Wgt_reg_542 <= Wgt_542;
		Wgt_reg_543 <= Wgt_543;
		Wgt_reg_544 <= Wgt_544;
		Wgt_reg_545 <= Wgt_545;
		Wgt_reg_546 <= Wgt_546;
		Wgt_reg_547 <= Wgt_547;
		Wgt_reg_548 <= Wgt_548;
		Wgt_reg_549 <= Wgt_549;
		Wgt_reg_550 <= Wgt_550;
		Wgt_reg_551 <= Wgt_551;
		Wgt_reg_552 <= Wgt_552;
		Wgt_reg_553 <= Wgt_553;
		Wgt_reg_554 <= Wgt_554;
		Wgt_reg_555 <= Wgt_555;
		Wgt_reg_556 <= Wgt_556;
		Wgt_reg_557 <= Wgt_557;
		Wgt_reg_558 <= Wgt_558;
		Wgt_reg_559 <= Wgt_559;
		Wgt_reg_560 <= Wgt_560;
		Wgt_reg_561 <= Wgt_561;
		Wgt_reg_562 <= Wgt_562;
		Wgt_reg_563 <= Wgt_563;
		Wgt_reg_564 <= Wgt_564;
		Wgt_reg_565 <= Wgt_565;
		Wgt_reg_566 <= Wgt_566;
		Wgt_reg_567 <= Wgt_567;
		Wgt_reg_568 <= Wgt_568;
		Wgt_reg_569 <= Wgt_569;
		Wgt_reg_570 <= Wgt_570;
		Wgt_reg_571 <= Wgt_571;
		Wgt_reg_572 <= Wgt_572;
		Wgt_reg_573 <= Wgt_573;
		Wgt_reg_574 <= Wgt_574;
		Wgt_reg_575 <= Wgt_575;
		Wgt_reg_576 <= Wgt_576;
		Wgt_reg_577 <= Wgt_577;
		Wgt_reg_578 <= Wgt_578;
		Wgt_reg_579 <= Wgt_579;
		Wgt_reg_580 <= Wgt_580;
		Wgt_reg_581 <= Wgt_581;
		Wgt_reg_582 <= Wgt_582;
		Wgt_reg_583 <= Wgt_583;
		Wgt_reg_584 <= Wgt_584;
		Wgt_reg_585 <= Wgt_585;
		Wgt_reg_586 <= Wgt_586;
		Wgt_reg_587 <= Wgt_587;
		Wgt_reg_588 <= Wgt_588;
		Wgt_reg_589 <= Wgt_589;
		Wgt_reg_590 <= Wgt_590;
		Wgt_reg_591 <= Wgt_591;
		Wgt_reg_592 <= Wgt_592;
		Wgt_reg_593 <= Wgt_593;
		Wgt_reg_594 <= Wgt_594;
		Wgt_reg_595 <= Wgt_595;
		Wgt_reg_596 <= Wgt_596;
		Wgt_reg_597 <= Wgt_597;
		Wgt_reg_598 <= Wgt_598;
		Wgt_reg_599 <= Wgt_599;
		Wgt_reg_600 <= Wgt_600;
		Wgt_reg_601 <= Wgt_601;
		Wgt_reg_602 <= Wgt_602;
		Wgt_reg_603 <= Wgt_603;
		Wgt_reg_604 <= Wgt_604;
		Wgt_reg_605 <= Wgt_605;
		Wgt_reg_606 <= Wgt_606;
		Wgt_reg_607 <= Wgt_607;
		Wgt_reg_608 <= Wgt_608;
		Wgt_reg_609 <= Wgt_609;
		Wgt_reg_610 <= Wgt_610;
		Wgt_reg_611 <= Wgt_611;
		Wgt_reg_612 <= Wgt_612;
		Wgt_reg_613 <= Wgt_613;
		Wgt_reg_614 <= Wgt_614;
		Wgt_reg_615 <= Wgt_615;
		Wgt_reg_616 <= Wgt_616;
		Wgt_reg_617 <= Wgt_617;
		Wgt_reg_618 <= Wgt_618;
		Wgt_reg_619 <= Wgt_619;
		Wgt_reg_620 <= Wgt_620;
		Wgt_reg_621 <= Wgt_621;
		Wgt_reg_622 <= Wgt_622;
		Wgt_reg_623 <= Wgt_623;
		Wgt_reg_624 <= Wgt_624;
		Wgt_reg_625 <= Wgt_625;
		Wgt_reg_626 <= Wgt_626;
		Wgt_reg_627 <= Wgt_627;
		Wgt_reg_628 <= Wgt_628;
		Wgt_reg_629 <= Wgt_629;
		Wgt_reg_630 <= Wgt_630;
		Wgt_reg_631 <= Wgt_631;
		Wgt_reg_632 <= Wgt_632;
		Wgt_reg_633 <= Wgt_633;
		Wgt_reg_634 <= Wgt_634;
		Wgt_reg_635 <= Wgt_635;
		Wgt_reg_636 <= Wgt_636;
		Wgt_reg_637 <= Wgt_637;
		Wgt_reg_638 <= Wgt_638;
		Wgt_reg_639 <= Wgt_639;
		Wgt_reg_640 <= Wgt_640;
		Wgt_reg_641 <= Wgt_641;
		Wgt_reg_642 <= Wgt_642;
		Wgt_reg_643 <= Wgt_643;
		Wgt_reg_644 <= Wgt_644;
		Wgt_reg_645 <= Wgt_645;
		Wgt_reg_646 <= Wgt_646;
		Wgt_reg_647 <= Wgt_647;
		Wgt_reg_648 <= Wgt_648;
		Wgt_reg_649 <= Wgt_649;
		Wgt_reg_650 <= Wgt_650;
		Wgt_reg_651 <= Wgt_651;
		Wgt_reg_652 <= Wgt_652;
		Wgt_reg_653 <= Wgt_653;
		Wgt_reg_654 <= Wgt_654;
		Wgt_reg_655 <= Wgt_655;
		Wgt_reg_656 <= Wgt_656;
		Wgt_reg_657 <= Wgt_657;
		Wgt_reg_658 <= Wgt_658;
		Wgt_reg_659 <= Wgt_659;
		Wgt_reg_660 <= Wgt_660;
		Wgt_reg_661 <= Wgt_661;
		Wgt_reg_662 <= Wgt_662;
		Wgt_reg_663 <= Wgt_663;
		Wgt_reg_664 <= Wgt_664;
		Wgt_reg_665 <= Wgt_665;
		Wgt_reg_666 <= Wgt_666;
		Wgt_reg_667 <= Wgt_667;
		Wgt_reg_668 <= Wgt_668;
		Wgt_reg_669 <= Wgt_669;
		Wgt_reg_670 <= Wgt_670;
		Wgt_reg_671 <= Wgt_671;
		Wgt_reg_672 <= Wgt_672;
		Wgt_reg_673 <= Wgt_673;
		Wgt_reg_674 <= Wgt_674;
		Wgt_reg_675 <= Wgt_675;
		Wgt_reg_676 <= Wgt_676;
		Wgt_reg_677 <= Wgt_677;
		Wgt_reg_678 <= Wgt_678;
		Wgt_reg_679 <= Wgt_679;
		Wgt_reg_680 <= Wgt_680;
		Wgt_reg_681 <= Wgt_681;
		Wgt_reg_682 <= Wgt_682;
		Wgt_reg_683 <= Wgt_683;
		Wgt_reg_684 <= Wgt_684;
		Wgt_reg_685 <= Wgt_685;
		Wgt_reg_686 <= Wgt_686;
		Wgt_reg_687 <= Wgt_687;
		Wgt_reg_688 <= Wgt_688;
		Wgt_reg_689 <= Wgt_689;
		Wgt_reg_690 <= Wgt_690;
		Wgt_reg_691 <= Wgt_691;
		Wgt_reg_692 <= Wgt_692;
		Wgt_reg_693 <= Wgt_693;
		Wgt_reg_694 <= Wgt_694;
		Wgt_reg_695 <= Wgt_695;
		Wgt_reg_696 <= Wgt_696;
		Wgt_reg_697 <= Wgt_697;
		Wgt_reg_698 <= Wgt_698;
		Wgt_reg_699 <= Wgt_699;
		Wgt_reg_700 <= Wgt_700;
		Wgt_reg_701 <= Wgt_701;
		Wgt_reg_702 <= Wgt_702;
		Wgt_reg_703 <= Wgt_703;
		Wgt_reg_704 <= Wgt_704;
		Wgt_reg_705 <= Wgt_705;
		Wgt_reg_706 <= Wgt_706;
		Wgt_reg_707 <= Wgt_707;
		Wgt_reg_708 <= Wgt_708;
		Wgt_reg_709 <= Wgt_709;
		Wgt_reg_710 <= Wgt_710;
		Wgt_reg_711 <= Wgt_711;
		Wgt_reg_712 <= Wgt_712;
		Wgt_reg_713 <= Wgt_713;
		Wgt_reg_714 <= Wgt_714;
		Wgt_reg_715 <= Wgt_715;
		Wgt_reg_716 <= Wgt_716;
		Wgt_reg_717 <= Wgt_717;
		Wgt_reg_718 <= Wgt_718;
		Wgt_reg_719 <= Wgt_719;
		Wgt_reg_720 <= Wgt_720;
		Wgt_reg_721 <= Wgt_721;
		Wgt_reg_722 <= Wgt_722;
		Wgt_reg_723 <= Wgt_723;
		Wgt_reg_724 <= Wgt_724;
		Wgt_reg_725 <= Wgt_725;
		Wgt_reg_726 <= Wgt_726;
		Wgt_reg_727 <= Wgt_727;
		Wgt_reg_728 <= Wgt_728;
		Wgt_reg_729 <= Wgt_729;
		Wgt_reg_730 <= Wgt_730;
		Wgt_reg_731 <= Wgt_731;
		Wgt_reg_732 <= Wgt_732;
		Wgt_reg_733 <= Wgt_733;
		Wgt_reg_734 <= Wgt_734;
		Wgt_reg_735 <= Wgt_735;
		Wgt_reg_736 <= Wgt_736;
		Wgt_reg_737 <= Wgt_737;
		Wgt_reg_738 <= Wgt_738;
		Wgt_reg_739 <= Wgt_739;
		Wgt_reg_740 <= Wgt_740;
		Wgt_reg_741 <= Wgt_741;
		Wgt_reg_742 <= Wgt_742;
		Wgt_reg_743 <= Wgt_743;
		Wgt_reg_744 <= Wgt_744;
		Wgt_reg_745 <= Wgt_745;
		Wgt_reg_746 <= Wgt_746;
		Wgt_reg_747 <= Wgt_747;
		Wgt_reg_748 <= Wgt_748;
		Wgt_reg_749 <= Wgt_749;
		Wgt_reg_750 <= Wgt_750;
		Wgt_reg_751 <= Wgt_751;
		Wgt_reg_752 <= Wgt_752;
		Wgt_reg_753 <= Wgt_753;
		Wgt_reg_754 <= Wgt_754;
		Wgt_reg_755 <= Wgt_755;
		Wgt_reg_756 <= Wgt_756;
		Wgt_reg_757 <= Wgt_757;
		Wgt_reg_758 <= Wgt_758;
		Wgt_reg_759 <= Wgt_759;
		Wgt_reg_760 <= Wgt_760;
		Wgt_reg_761 <= Wgt_761;
		Wgt_reg_762 <= Wgt_762;
		Wgt_reg_763 <= Wgt_763;
		Wgt_reg_764 <= Wgt_764;
		Wgt_reg_765 <= Wgt_765;
		Wgt_reg_766 <= Wgt_766;
		Wgt_reg_767 <= Wgt_767;
		Wgt_reg_768 <= Wgt_768;
		Wgt_reg_769 <= Wgt_769;
		Wgt_reg_770 <= Wgt_770;
		Wgt_reg_771 <= Wgt_771;
		Wgt_reg_772 <= Wgt_772;
		Wgt_reg_773 <= Wgt_773;
		Wgt_reg_774 <= Wgt_774;
		Wgt_reg_775 <= Wgt_775;
		Wgt_reg_776 <= Wgt_776;
		Wgt_reg_777 <= Wgt_777;
		Wgt_reg_778 <= Wgt_778;
		Wgt_reg_779 <= Wgt_779;
		Wgt_reg_780 <= Wgt_780;
		Wgt_reg_781 <= Wgt_781;
		Wgt_reg_782 <= Wgt_782;
		Wgt_reg_783 <= Wgt_783;
		Wgt_reg_784 <= Wgt_784;

			
			state<=48;
			end
			else begin state<= 7'b0000000; end
		end

		48: begin
			select <= 6'b000000;
			state <= 7'b0000001; 
		end

		7'b0000001: begin
			select<=6'b000001;
			state<=7'b0000010;
		end
		7'b0000010: begin
			select<=2;
			state<=3;
		end
		3: begin
			select<=3;
			state<=4;
		end
		4:begin
			select<=4;
			state<=5;
		end
		5:begin
			select<=5;
			state<=6;
		end
		6:begin  //1st mul???
			select<=6;
			state<=7;
		end
		7: begin  //1st mul
			select<=7;
			state<=8;
		end
		8: begin
			select<=8;
			state<=9;
		end
		9: begin
			select<=9;
			state<=10;
		end
		10: begin
			select<=10;
			state<=11;
		end
		11:begin
			select<=11;
			state<=12;
		end
		12:begin
			select<=12;
			state<=13;
		end
		13:begin
			select<=13;
			state<=14;
		end
		14: begin
			select<=14;
			state<=15;
		end
		15: begin
			select<=15;
			state<=16;
		end
		16: begin
			select<=16;
			//sum_reg0<=sum;
			state<=17;
		end
		17: begin
			select<=17;
			sum_reg0<=sum;
			state<=18;
		end
		18:begin
			select<=18;
			sum_reg1<=sum;
			state<=19;
		end
		19:begin
			select<=19;
			sum_reg2<=sum;
			state<=20;
			
		end
		20:begin
			select<=20;
			sum_reg3<=sum;
			state<=21;

		end
		21:begin
			select<=21;
			sum_reg4<=sum;
			state<=22;
		end
		22:begin
			select<=22;
			sum_reg5<=sum;
			state<=23;
		end
		23: begin
			select<=23;
			sum_reg6<=sum;
			state<=24;
		end
		24: begin
			select<=24;
			sum_reg7<=sum;
			state<=25;
		end
		25: begin
			select<=25;
			sum_reg8<=sum;
			state<=26;
		end
		26: begin
			select<=26;
			sum_reg9<=sum;
			state<=27;
		end
		27:begin
			select<=27;
			sum_reg10<=sum;
			state<=28;
		end
		28:begin
			sum_reg11<=sum;
			state<=29;
		end
		29:begin
		sum_reg12<=sum;
		state<=30;
		end

		30:begin
		sum_reg13<=sum;
		state<=31;
		end

		31:begin
		sum_reg14<=sum;
		state<=32;
		end

		32:begin
		sum_reg15<=sum;
		state<=33;
		end

		33:begin
		sum_reg16<=sum;
		state<=34;
		end

		34:begin
		sum_reg17<=sum;
		state<=35;
		end

		35:begin
		sum_reg18<=sum;
		state<=36;
		end

		36:begin
		sum_reg19<=sum;
		state<=37;
		end

		37:begin
		sum_reg20<=sum;
		state<=38;
		end

		38:begin
		sum_reg21<=sum;
		state<=39;
		end

		39:begin
		sum_reg22<=sum;
		state<=40;
		end

		40:begin
		sum_reg23<=sum;
		state<=41;
		end

		41:begin
		sum_reg24<=sum;
		state<=42;
		end

		42:begin
		sum_reg25<=sum;
		state<=43;
		end

		43:begin
		sum_reg26<=sum;
		state<=44;
		end

		44:begin
		sum_reg27<=sum;
		state<= 45;//7'b0000000;
		end

		45:begin
			  sum_sim_reg0<=sum_reg0;
			  sum_sim_reg1<=sum_reg1;
			  sum_sim_reg2<=sum_reg2;
			  sum_sim_reg3<=sum_reg3;
			  sum_sim_reg4<=sum_reg4;
			  sum_sim_reg5<=sum_reg5;
			  sum_sim_reg6<=sum_reg6;
			  sum_sim_reg7<=sum_reg7;
			  sum_sim_reg8<=sum_reg8;
			  sum_sim_reg9<=sum_reg9;
			  sum_sim_reg10<=sum_reg10;
			  sum_sim_reg11<=sum_reg11;
			  sum_sim_reg12<=sum_reg12;
			  sum_sim_reg13<=sum_reg13;
			  sum_sim_reg14<=sum_reg14;
			  sum_sim_reg15<=sum_reg15;
			  sum_sim_reg16<=sum_reg16;
			  sum_sim_reg17<=sum_reg17;
			  sum_sim_reg18<=sum_reg18;
			  sum_sim_reg19<=sum_reg19;
			  sum_sim_reg20<=sum_reg20;
			  sum_sim_reg21<=sum_reg21;
			  sum_sim_reg22<=sum_reg22;
			  sum_sim_reg23<=sum_reg23;
			  sum_sim_reg24<=sum_reg24;
			  sum_sim_reg25<=sum_reg25;
			  sum_sim_reg26<=sum_reg26;
			  sum_sim_reg27<=sum_reg27;
			  counter<=0;
			  state <=46;
		end
		46: begin
			state<=(counter<23)?46:47; //大概转50多次确保算完sum
			counter<=counter+1;
		end
		47: begin
			cell_out_r <= tot_out_real;
			Output_Valid_r <= 1'b1;
			state <= 7'b0000000;
		end
		default:begin
			
			state<=7'b0000000; 
		end


	endcase

	end
end

assign cell_out = cell_out_r;
assign Output_Valid = Output_Valid_r;
endmodule
